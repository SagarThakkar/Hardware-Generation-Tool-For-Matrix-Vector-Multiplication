include "s_thakkar_mvm_4_4_8_1.sv";
// Testbench, with parameters k=4, p=4, b=8, g=1

//This Test bench shows values on normal computation and in the next cycle only the vector is updated keeping the matrix same
 module tb1();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb1");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadVector=1;
@(posedge clk);
#1; loadVector=0;
data_in = 1;
@(posedge clk);
#1;data_in = -3;
@(posedge clk);
#1;data_in = -4;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
//This testbench incorporates two iterations in the first iteration the values are computed according to the values and in the next iteration only the Matrix is updated keeping vector
module tb2();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

// Set input values.
initial begin  
start = 0; reset = 1;data_in=8'bx;
@(posedge clk);
#1; reset=0;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge clk);
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
start=0; reset=1; data_in=8'bx;
@(posedge clk);
#1; reset=0; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0; data_in = 1;
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
#1;data_in = 5;
@(posedge clk);
#1;data_in = 6;
@(posedge clk);
#1;data_in = 7;
@(posedge clk);
#1;data_in = 8;
@(posedge clk);
#1;data_in = 9;
@(posedge clk);
#1;data_in = 10;
@(posedge clk);
#1;data_in = 11;
@(posedge clk);
#1;data_in = 12;
@(posedge clk);
#1;data_in = 13;
@(posedge clk);
#1;data_in = 14;
@(posedge clk);
#1;data_in = 15;
@(posedge clk);
#1;data_in = 16;
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=1; 
@(posedge clk);
#1;data_in = 2;
@(posedge clk);
#1;data_in = 3;
@(posedge clk);
#1;data_in = 4;
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

integer filehandle=$fopen("proj3_outValuestb2");
// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; loadMatrix=1;
@(posedge clk);
#1; loadMatrix=0;
data_in = 1;
@(posedge clk);
#1;data_in = -5;
@(posedge clk);
#1;data_in = -6;
@(posedge clk);
#1;data_in = -7;
@(posedge clk);
#1;data_in = -8;
@(posedge clk);
#1;data_in = -9;
@(posedge clk);
#1;data_in = -10;
@(posedge clk);
#1;data_in = -11;
@(posedge clk);
#1;data_in = -12;
@(posedge clk);
#1;data_in = -13;
@(posedge clk);
#1;data_in = -14;
@(posedge clk);
#1;data_in = -15;
@(posedge clk);
#1;data_in = -16;
@(posedge clk);
#1;data_in = -17;
@(posedge clk);
#1;data_in = -18;
@(posedge clk);
#1;data_in = -19;
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=4, p=4, b=8, g=1

module tb3();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData3[19:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb3", testData3);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb3");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData3[0];
@(posedge clk);
#1;data_in = testData3[1];
@(posedge clk);
#1;data_in = testData3[2];
@(posedge clk);
#1;data_in = testData3[3];
@(posedge clk);
#1;data_in = testData3[4];
@(posedge clk);
#1;data_in = testData3[5];
@(posedge clk);
#1;data_in = testData3[6];
@(posedge clk);
#1;data_in = testData3[7];
@(posedge clk);
#1;data_in = testData3[8];
@(posedge clk);
#1;data_in = testData3[9];
@(posedge clk);
#1;data_in = testData3[10];
@(posedge clk);
#1;data_in = testData3[11];
@(posedge clk);
#1;data_in = testData3[12];
@(posedge clk);
#1;data_in = testData3[13];
@(posedge clk);
#1;data_in = testData3[14];
@(posedge clk);
#1;data_in = testData3[15];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData3[16]; 
@(posedge clk);
#1;data_in = testData3[17];
@(posedge clk);
#1;data_in = testData3[18];
@(posedge clk);
#1;data_in = testData3[19];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=4, p=4, b=8, g=1

module tb4();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData4[219:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb4", testData4);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb4");
  initial begin 
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData4[0];
@(posedge clk);
#1;data_in = testData4[1];
@(posedge clk);
#1;data_in = testData4[2];
@(posedge clk);
#1;data_in = testData4[3];
@(posedge clk);
#1;data_in = testData4[4];
@(posedge clk);
#1;data_in = testData4[5];
@(posedge clk);
#1;data_in = testData4[6];
@(posedge clk);
#1;data_in = testData4[7];
@(posedge clk);
#1;data_in = testData4[8];
@(posedge clk);
#1;data_in = testData4[9];
@(posedge clk);
#1;data_in = testData4[10];
@(posedge clk);
#1;data_in = testData4[11];
@(posedge clk);
#1;data_in = testData4[12];
@(posedge clk);
#1;data_in = testData4[13];
@(posedge clk);
#1;data_in = testData4[14];
@(posedge clk);
#1;data_in = testData4[15];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData4[16]; 
@(posedge clk);
#1;data_in = testData4[17];
@(posedge clk);
#1;data_in = testData4[18];
@(posedge clk);
#1;data_in = testData4[19];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 end

// wait for done signal and output  
initial begin
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[20]; 
@(posedge clk);
#1;data_in = testData4[21];
@(posedge clk);
#1;data_in = testData4[22];
@(posedge clk);
#1;data_in = testData4[23];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[24]; 
@(posedge clk);
#1;data_in = testData4[25];
@(posedge clk);
#1;data_in = testData4[26];
@(posedge clk);
#1;data_in = testData4[27];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[28]; 
@(posedge clk);
#1;data_in = testData4[29];
@(posedge clk);
#1;data_in = testData4[30];
@(posedge clk);
#1;data_in = testData4[31];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[32]; 
@(posedge clk);
#1;data_in = testData4[33];
@(posedge clk);
#1;data_in = testData4[34];
@(posedge clk);
#1;data_in = testData4[35];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[36]; 
@(posedge clk);
#1;data_in = testData4[37];
@(posedge clk);
#1;data_in = testData4[38];
@(posedge clk);
#1;data_in = testData4[39];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[40]; 
@(posedge clk);
#1;data_in = testData4[41];
@(posedge clk);
#1;data_in = testData4[42];
@(posedge clk);
#1;data_in = testData4[43];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[44]; 
@(posedge clk);
#1;data_in = testData4[45];
@(posedge clk);
#1;data_in = testData4[46];
@(posedge clk);
#1;data_in = testData4[47];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[48]; 
@(posedge clk);
#1;data_in = testData4[49];
@(posedge clk);
#1;data_in = testData4[50];
@(posedge clk);
#1;data_in = testData4[51];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[52]; 
@(posedge clk);
#1;data_in = testData4[53];
@(posedge clk);
#1;data_in = testData4[54];
@(posedge clk);
#1;data_in = testData4[55];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[56]; 
@(posedge clk);
#1;data_in = testData4[57];
@(posedge clk);
#1;data_in = testData4[58];
@(posedge clk);
#1;data_in = testData4[59];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[60]; 
@(posedge clk);
#1;data_in = testData4[61];
@(posedge clk);
#1;data_in = testData4[62];
@(posedge clk);
#1;data_in = testData4[63];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[64]; 
@(posedge clk);
#1;data_in = testData4[65];
@(posedge clk);
#1;data_in = testData4[66];
@(posedge clk);
#1;data_in = testData4[67];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[68]; 
@(posedge clk);
#1;data_in = testData4[69];
@(posedge clk);
#1;data_in = testData4[70];
@(posedge clk);
#1;data_in = testData4[71];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[72]; 
@(posedge clk);
#1;data_in = testData4[73];
@(posedge clk);
#1;data_in = testData4[74];
@(posedge clk);
#1;data_in = testData4[75];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[76]; 
@(posedge clk);
#1;data_in = testData4[77];
@(posedge clk);
#1;data_in = testData4[78];
@(posedge clk);
#1;data_in = testData4[79];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[80]; 
@(posedge clk);
#1;data_in = testData4[81];
@(posedge clk);
#1;data_in = testData4[82];
@(posedge clk);
#1;data_in = testData4[83];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[84]; 
@(posedge clk);
#1;data_in = testData4[85];
@(posedge clk);
#1;data_in = testData4[86];
@(posedge clk);
#1;data_in = testData4[87];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[88]; 
@(posedge clk);
#1;data_in = testData4[89];
@(posedge clk);
#1;data_in = testData4[90];
@(posedge clk);
#1;data_in = testData4[91];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[92]; 
@(posedge clk);
#1;data_in = testData4[93];
@(posedge clk);
#1;data_in = testData4[94];
@(posedge clk);
#1;data_in = testData4[95];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[96]; 
@(posedge clk);
#1;data_in = testData4[97];
@(posedge clk);
#1;data_in = testData4[98];
@(posedge clk);
#1;data_in = testData4[99];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[100]; 
@(posedge clk);
#1;data_in = testData4[101];
@(posedge clk);
#1;data_in = testData4[102];
@(posedge clk);
#1;data_in = testData4[103];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[104]; 
@(posedge clk);
#1;data_in = testData4[105];
@(posedge clk);
#1;data_in = testData4[106];
@(posedge clk);
#1;data_in = testData4[107];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[108]; 
@(posedge clk);
#1;data_in = testData4[109];
@(posedge clk);
#1;data_in = testData4[110];
@(posedge clk);
#1;data_in = testData4[111];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[112]; 
@(posedge clk);
#1;data_in = testData4[113];
@(posedge clk);
#1;data_in = testData4[114];
@(posedge clk);
#1;data_in = testData4[115];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[116]; 
@(posedge clk);
#1;data_in = testData4[117];
@(posedge clk);
#1;data_in = testData4[118];
@(posedge clk);
#1;data_in = testData4[119];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[120]; 
@(posedge clk);
#1;data_in = testData4[121];
@(posedge clk);
#1;data_in = testData4[122];
@(posedge clk);
#1;data_in = testData4[123];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[124]; 
@(posedge clk);
#1;data_in = testData4[125];
@(posedge clk);
#1;data_in = testData4[126];
@(posedge clk);
#1;data_in = testData4[127];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[128]; 
@(posedge clk);
#1;data_in = testData4[129];
@(posedge clk);
#1;data_in = testData4[130];
@(posedge clk);
#1;data_in = testData4[131];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[132]; 
@(posedge clk);
#1;data_in = testData4[133];
@(posedge clk);
#1;data_in = testData4[134];
@(posedge clk);
#1;data_in = testData4[135];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[136]; 
@(posedge clk);
#1;data_in = testData4[137];
@(posedge clk);
#1;data_in = testData4[138];
@(posedge clk);
#1;data_in = testData4[139];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[140]; 
@(posedge clk);
#1;data_in = testData4[141];
@(posedge clk);
#1;data_in = testData4[142];
@(posedge clk);
#1;data_in = testData4[143];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[144]; 
@(posedge clk);
#1;data_in = testData4[145];
@(posedge clk);
#1;data_in = testData4[146];
@(posedge clk);
#1;data_in = testData4[147];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[148]; 
@(posedge clk);
#1;data_in = testData4[149];
@(posedge clk);
#1;data_in = testData4[150];
@(posedge clk);
#1;data_in = testData4[151];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[152]; 
@(posedge clk);
#1;data_in = testData4[153];
@(posedge clk);
#1;data_in = testData4[154];
@(posedge clk);
#1;data_in = testData4[155];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[156]; 
@(posedge clk);
#1;data_in = testData4[157];
@(posedge clk);
#1;data_in = testData4[158];
@(posedge clk);
#1;data_in = testData4[159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[160]; 
@(posedge clk);
#1;data_in = testData4[161];
@(posedge clk);
#1;data_in = testData4[162];
@(posedge clk);
#1;data_in = testData4[163];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[164]; 
@(posedge clk);
#1;data_in = testData4[165];
@(posedge clk);
#1;data_in = testData4[166];
@(posedge clk);
#1;data_in = testData4[167];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[168]; 
@(posedge clk);
#1;data_in = testData4[169];
@(posedge clk);
#1;data_in = testData4[170];
@(posedge clk);
#1;data_in = testData4[171];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[172]; 
@(posedge clk);
#1;data_in = testData4[173];
@(posedge clk);
#1;data_in = testData4[174];
@(posedge clk);
#1;data_in = testData4[175];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[176]; 
@(posedge clk);
#1;data_in = testData4[177];
@(posedge clk);
#1;data_in = testData4[178];
@(posedge clk);
#1;data_in = testData4[179];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[180]; 
@(posedge clk);
#1;data_in = testData4[181];
@(posedge clk);
#1;data_in = testData4[182];
@(posedge clk);
#1;data_in = testData4[183];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[184]; 
@(posedge clk);
#1;data_in = testData4[185];
@(posedge clk);
#1;data_in = testData4[186];
@(posedge clk);
#1;data_in = testData4[187];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[188]; 
@(posedge clk);
#1;data_in = testData4[189];
@(posedge clk);
#1;data_in = testData4[190];
@(posedge clk);
#1;data_in = testData4[191];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[192]; 
@(posedge clk);
#1;data_in = testData4[193];
@(posedge clk);
#1;data_in = testData4[194];
@(posedge clk);
#1;data_in = testData4[195];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[196]; 
@(posedge clk);
#1;data_in = testData4[197];
@(posedge clk);
#1;data_in = testData4[198];
@(posedge clk);
#1;data_in = testData4[199];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[200]; 
@(posedge clk);
#1;data_in = testData4[201];
@(posedge clk);
#1;data_in = testData4[202];
@(posedge clk);
#1;data_in = testData4[203];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[204]; 
@(posedge clk);
#1;data_in = testData4[205];
@(posedge clk);
#1;data_in = testData4[206];
@(posedge clk);
#1;data_in = testData4[207];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[208]; 
@(posedge clk);
#1;data_in = testData4[209];
@(posedge clk);
#1;data_in = testData4[210];
@(posedge clk);
#1;data_in = testData4[211];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[212]; 
@(posedge clk);
#1;data_in = testData4[213];
@(posedge clk);
#1;data_in = testData4[214];
@(posedge clk);
#1;data_in = testData4[215];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadVector =1;
@(posedge clk);
#1 ; loadVector =0;
data_in=testData4[216]; 
@(posedge clk);
#1;data_in = testData4[217];
@(posedge clk);
#1;data_in = testData4[218];
@(posedge clk);
#1;data_in = testData4[219];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
module tb6();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData6[1019:0];
   //read input from C file inputDatapart2     
 initial $readmemh("proj3_inputDatatb6", testData6);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb6");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[0];
@(posedge clk);
#1;data_in = testData6[1];
@(posedge clk);
#1;data_in = testData6[2];
@(posedge clk);
#1;data_in = testData6[3];
@(posedge clk);
#1;data_in = testData6[4];
@(posedge clk);
#1;data_in = testData6[5];
@(posedge clk);
#1;data_in = testData6[6];
@(posedge clk);
#1;data_in = testData6[7];
@(posedge clk);
#1;data_in = testData6[8];
@(posedge clk);
#1;data_in = testData6[9];
@(posedge clk);
#1;data_in = testData6[10];
@(posedge clk);
#1;data_in = testData6[11];
@(posedge clk);
#1;data_in = testData6[12];
@(posedge clk);
#1;data_in = testData6[13];
@(posedge clk);
#1;data_in = testData6[14];
@(posedge clk);
#1;data_in = testData6[15];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[16]; 
@(posedge clk);
#1;data_in = testData6[17];
@(posedge clk);
#1;data_in = testData6[18];
@(posedge clk);
#1;data_in = testData6[19];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[20];
@(posedge clk);
#1;data_in = testData6[21];
@(posedge clk);
#1;data_in = testData6[22];
@(posedge clk);
#1;data_in = testData6[23];
@(posedge clk);
#1;data_in = testData6[24];
@(posedge clk);
#1;data_in = testData6[25];
@(posedge clk);
#1;data_in = testData6[26];
@(posedge clk);
#1;data_in = testData6[27];
@(posedge clk);
#1;data_in = testData6[28];
@(posedge clk);
#1;data_in = testData6[29];
@(posedge clk);
#1;data_in = testData6[30];
@(posedge clk);
#1;data_in = testData6[31];
@(posedge clk);
#1;data_in = testData6[32];
@(posedge clk);
#1;data_in = testData6[33];
@(posedge clk);
#1;data_in = testData6[34];
@(posedge clk);
#1;data_in = testData6[35];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[36]; 
@(posedge clk);
#1;data_in = testData6[37];
@(posedge clk);
#1;data_in = testData6[38];
@(posedge clk);
#1;data_in = testData6[39];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[40];
@(posedge clk);
#1;data_in = testData6[41];
@(posedge clk);
#1;data_in = testData6[42];
@(posedge clk);
#1;data_in = testData6[43];
@(posedge clk);
#1;data_in = testData6[44];
@(posedge clk);
#1;data_in = testData6[45];
@(posedge clk);
#1;data_in = testData6[46];
@(posedge clk);
#1;data_in = testData6[47];
@(posedge clk);
#1;data_in = testData6[48];
@(posedge clk);
#1;data_in = testData6[49];
@(posedge clk);
#1;data_in = testData6[50];
@(posedge clk);
#1;data_in = testData6[51];
@(posedge clk);
#1;data_in = testData6[52];
@(posedge clk);
#1;data_in = testData6[53];
@(posedge clk);
#1;data_in = testData6[54];
@(posedge clk);
#1;data_in = testData6[55];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[56]; 
@(posedge clk);
#1;data_in = testData6[57];
@(posedge clk);
#1;data_in = testData6[58];
@(posedge clk);
#1;data_in = testData6[59];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[60];
@(posedge clk);
#1;data_in = testData6[61];
@(posedge clk);
#1;data_in = testData6[62];
@(posedge clk);
#1;data_in = testData6[63];
@(posedge clk);
#1;data_in = testData6[64];
@(posedge clk);
#1;data_in = testData6[65];
@(posedge clk);
#1;data_in = testData6[66];
@(posedge clk);
#1;data_in = testData6[67];
@(posedge clk);
#1;data_in = testData6[68];
@(posedge clk);
#1;data_in = testData6[69];
@(posedge clk);
#1;data_in = testData6[70];
@(posedge clk);
#1;data_in = testData6[71];
@(posedge clk);
#1;data_in = testData6[72];
@(posedge clk);
#1;data_in = testData6[73];
@(posedge clk);
#1;data_in = testData6[74];
@(posedge clk);
#1;data_in = testData6[75];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[76]; 
@(posedge clk);
#1;data_in = testData6[77];
@(posedge clk);
#1;data_in = testData6[78];
@(posedge clk);
#1;data_in = testData6[79];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[80];
@(posedge clk);
#1;data_in = testData6[81];
@(posedge clk);
#1;data_in = testData6[82];
@(posedge clk);
#1;data_in = testData6[83];
@(posedge clk);
#1;data_in = testData6[84];
@(posedge clk);
#1;data_in = testData6[85];
@(posedge clk);
#1;data_in = testData6[86];
@(posedge clk);
#1;data_in = testData6[87];
@(posedge clk);
#1;data_in = testData6[88];
@(posedge clk);
#1;data_in = testData6[89];
@(posedge clk);
#1;data_in = testData6[90];
@(posedge clk);
#1;data_in = testData6[91];
@(posedge clk);
#1;data_in = testData6[92];
@(posedge clk);
#1;data_in = testData6[93];
@(posedge clk);
#1;data_in = testData6[94];
@(posedge clk);
#1;data_in = testData6[95];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[96]; 
@(posedge clk);
#1;data_in = testData6[97];
@(posedge clk);
#1;data_in = testData6[98];
@(posedge clk);
#1;data_in = testData6[99];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[100];
@(posedge clk);
#1;data_in = testData6[101];
@(posedge clk);
#1;data_in = testData6[102];
@(posedge clk);
#1;data_in = testData6[103];
@(posedge clk);
#1;data_in = testData6[104];
@(posedge clk);
#1;data_in = testData6[105];
@(posedge clk);
#1;data_in = testData6[106];
@(posedge clk);
#1;data_in = testData6[107];
@(posedge clk);
#1;data_in = testData6[108];
@(posedge clk);
#1;data_in = testData6[109];
@(posedge clk);
#1;data_in = testData6[110];
@(posedge clk);
#1;data_in = testData6[111];
@(posedge clk);
#1;data_in = testData6[112];
@(posedge clk);
#1;data_in = testData6[113];
@(posedge clk);
#1;data_in = testData6[114];
@(posedge clk);
#1;data_in = testData6[115];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[116]; 
@(posedge clk);
#1;data_in = testData6[117];
@(posedge clk);
#1;data_in = testData6[118];
@(posedge clk);
#1;data_in = testData6[119];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[120];
@(posedge clk);
#1;data_in = testData6[121];
@(posedge clk);
#1;data_in = testData6[122];
@(posedge clk);
#1;data_in = testData6[123];
@(posedge clk);
#1;data_in = testData6[124];
@(posedge clk);
#1;data_in = testData6[125];
@(posedge clk);
#1;data_in = testData6[126];
@(posedge clk);
#1;data_in = testData6[127];
@(posedge clk);
#1;data_in = testData6[128];
@(posedge clk);
#1;data_in = testData6[129];
@(posedge clk);
#1;data_in = testData6[130];
@(posedge clk);
#1;data_in = testData6[131];
@(posedge clk);
#1;data_in = testData6[132];
@(posedge clk);
#1;data_in = testData6[133];
@(posedge clk);
#1;data_in = testData6[134];
@(posedge clk);
#1;data_in = testData6[135];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[136]; 
@(posedge clk);
#1;data_in = testData6[137];
@(posedge clk);
#1;data_in = testData6[138];
@(posedge clk);
#1;data_in = testData6[139];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[140];
@(posedge clk);
#1;data_in = testData6[141];
@(posedge clk);
#1;data_in = testData6[142];
@(posedge clk);
#1;data_in = testData6[143];
@(posedge clk);
#1;data_in = testData6[144];
@(posedge clk);
#1;data_in = testData6[145];
@(posedge clk);
#1;data_in = testData6[146];
@(posedge clk);
#1;data_in = testData6[147];
@(posedge clk);
#1;data_in = testData6[148];
@(posedge clk);
#1;data_in = testData6[149];
@(posedge clk);
#1;data_in = testData6[150];
@(posedge clk);
#1;data_in = testData6[151];
@(posedge clk);
#1;data_in = testData6[152];
@(posedge clk);
#1;data_in = testData6[153];
@(posedge clk);
#1;data_in = testData6[154];
@(posedge clk);
#1;data_in = testData6[155];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[156]; 
@(posedge clk);
#1;data_in = testData6[157];
@(posedge clk);
#1;data_in = testData6[158];
@(posedge clk);
#1;data_in = testData6[159];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[160];
@(posedge clk);
#1;data_in = testData6[161];
@(posedge clk);
#1;data_in = testData6[162];
@(posedge clk);
#1;data_in = testData6[163];
@(posedge clk);
#1;data_in = testData6[164];
@(posedge clk);
#1;data_in = testData6[165];
@(posedge clk);
#1;data_in = testData6[166];
@(posedge clk);
#1;data_in = testData6[167];
@(posedge clk);
#1;data_in = testData6[168];
@(posedge clk);
#1;data_in = testData6[169];
@(posedge clk);
#1;data_in = testData6[170];
@(posedge clk);
#1;data_in = testData6[171];
@(posedge clk);
#1;data_in = testData6[172];
@(posedge clk);
#1;data_in = testData6[173];
@(posedge clk);
#1;data_in = testData6[174];
@(posedge clk);
#1;data_in = testData6[175];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[176]; 
@(posedge clk);
#1;data_in = testData6[177];
@(posedge clk);
#1;data_in = testData6[178];
@(posedge clk);
#1;data_in = testData6[179];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[180];
@(posedge clk);
#1;data_in = testData6[181];
@(posedge clk);
#1;data_in = testData6[182];
@(posedge clk);
#1;data_in = testData6[183];
@(posedge clk);
#1;data_in = testData6[184];
@(posedge clk);
#1;data_in = testData6[185];
@(posedge clk);
#1;data_in = testData6[186];
@(posedge clk);
#1;data_in = testData6[187];
@(posedge clk);
#1;data_in = testData6[188];
@(posedge clk);
#1;data_in = testData6[189];
@(posedge clk);
#1;data_in = testData6[190];
@(posedge clk);
#1;data_in = testData6[191];
@(posedge clk);
#1;data_in = testData6[192];
@(posedge clk);
#1;data_in = testData6[193];
@(posedge clk);
#1;data_in = testData6[194];
@(posedge clk);
#1;data_in = testData6[195];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[196]; 
@(posedge clk);
#1;data_in = testData6[197];
@(posedge clk);
#1;data_in = testData6[198];
@(posedge clk);
#1;data_in = testData6[199];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[200];
@(posedge clk);
#1;data_in = testData6[201];
@(posedge clk);
#1;data_in = testData6[202];
@(posedge clk);
#1;data_in = testData6[203];
@(posedge clk);
#1;data_in = testData6[204];
@(posedge clk);
#1;data_in = testData6[205];
@(posedge clk);
#1;data_in = testData6[206];
@(posedge clk);
#1;data_in = testData6[207];
@(posedge clk);
#1;data_in = testData6[208];
@(posedge clk);
#1;data_in = testData6[209];
@(posedge clk);
#1;data_in = testData6[210];
@(posedge clk);
#1;data_in = testData6[211];
@(posedge clk);
#1;data_in = testData6[212];
@(posedge clk);
#1;data_in = testData6[213];
@(posedge clk);
#1;data_in = testData6[214];
@(posedge clk);
#1;data_in = testData6[215];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[216]; 
@(posedge clk);
#1;data_in = testData6[217];
@(posedge clk);
#1;data_in = testData6[218];
@(posedge clk);
#1;data_in = testData6[219];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[220];
@(posedge clk);
#1;data_in = testData6[221];
@(posedge clk);
#1;data_in = testData6[222];
@(posedge clk);
#1;data_in = testData6[223];
@(posedge clk);
#1;data_in = testData6[224];
@(posedge clk);
#1;data_in = testData6[225];
@(posedge clk);
#1;data_in = testData6[226];
@(posedge clk);
#1;data_in = testData6[227];
@(posedge clk);
#1;data_in = testData6[228];
@(posedge clk);
#1;data_in = testData6[229];
@(posedge clk);
#1;data_in = testData6[230];
@(posedge clk);
#1;data_in = testData6[231];
@(posedge clk);
#1;data_in = testData6[232];
@(posedge clk);
#1;data_in = testData6[233];
@(posedge clk);
#1;data_in = testData6[234];
@(posedge clk);
#1;data_in = testData6[235];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[236]; 
@(posedge clk);
#1;data_in = testData6[237];
@(posedge clk);
#1;data_in = testData6[238];
@(posedge clk);
#1;data_in = testData6[239];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[240];
@(posedge clk);
#1;data_in = testData6[241];
@(posedge clk);
#1;data_in = testData6[242];
@(posedge clk);
#1;data_in = testData6[243];
@(posedge clk);
#1;data_in = testData6[244];
@(posedge clk);
#1;data_in = testData6[245];
@(posedge clk);
#1;data_in = testData6[246];
@(posedge clk);
#1;data_in = testData6[247];
@(posedge clk);
#1;data_in = testData6[248];
@(posedge clk);
#1;data_in = testData6[249];
@(posedge clk);
#1;data_in = testData6[250];
@(posedge clk);
#1;data_in = testData6[251];
@(posedge clk);
#1;data_in = testData6[252];
@(posedge clk);
#1;data_in = testData6[253];
@(posedge clk);
#1;data_in = testData6[254];
@(posedge clk);
#1;data_in = testData6[255];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[256]; 
@(posedge clk);
#1;data_in = testData6[257];
@(posedge clk);
#1;data_in = testData6[258];
@(posedge clk);
#1;data_in = testData6[259];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[260];
@(posedge clk);
#1;data_in = testData6[261];
@(posedge clk);
#1;data_in = testData6[262];
@(posedge clk);
#1;data_in = testData6[263];
@(posedge clk);
#1;data_in = testData6[264];
@(posedge clk);
#1;data_in = testData6[265];
@(posedge clk);
#1;data_in = testData6[266];
@(posedge clk);
#1;data_in = testData6[267];
@(posedge clk);
#1;data_in = testData6[268];
@(posedge clk);
#1;data_in = testData6[269];
@(posedge clk);
#1;data_in = testData6[270];
@(posedge clk);
#1;data_in = testData6[271];
@(posedge clk);
#1;data_in = testData6[272];
@(posedge clk);
#1;data_in = testData6[273];
@(posedge clk);
#1;data_in = testData6[274];
@(posedge clk);
#1;data_in = testData6[275];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[276]; 
@(posedge clk);
#1;data_in = testData6[277];
@(posedge clk);
#1;data_in = testData6[278];
@(posedge clk);
#1;data_in = testData6[279];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[280];
@(posedge clk);
#1;data_in = testData6[281];
@(posedge clk);
#1;data_in = testData6[282];
@(posedge clk);
#1;data_in = testData6[283];
@(posedge clk);
#1;data_in = testData6[284];
@(posedge clk);
#1;data_in = testData6[285];
@(posedge clk);
#1;data_in = testData6[286];
@(posedge clk);
#1;data_in = testData6[287];
@(posedge clk);
#1;data_in = testData6[288];
@(posedge clk);
#1;data_in = testData6[289];
@(posedge clk);
#1;data_in = testData6[290];
@(posedge clk);
#1;data_in = testData6[291];
@(posedge clk);
#1;data_in = testData6[292];
@(posedge clk);
#1;data_in = testData6[293];
@(posedge clk);
#1;data_in = testData6[294];
@(posedge clk);
#1;data_in = testData6[295];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[296]; 
@(posedge clk);
#1;data_in = testData6[297];
@(posedge clk);
#1;data_in = testData6[298];
@(posedge clk);
#1;data_in = testData6[299];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[300];
@(posedge clk);
#1;data_in = testData6[301];
@(posedge clk);
#1;data_in = testData6[302];
@(posedge clk);
#1;data_in = testData6[303];
@(posedge clk);
#1;data_in = testData6[304];
@(posedge clk);
#1;data_in = testData6[305];
@(posedge clk);
#1;data_in = testData6[306];
@(posedge clk);
#1;data_in = testData6[307];
@(posedge clk);
#1;data_in = testData6[308];
@(posedge clk);
#1;data_in = testData6[309];
@(posedge clk);
#1;data_in = testData6[310];
@(posedge clk);
#1;data_in = testData6[311];
@(posedge clk);
#1;data_in = testData6[312];
@(posedge clk);
#1;data_in = testData6[313];
@(posedge clk);
#1;data_in = testData6[314];
@(posedge clk);
#1;data_in = testData6[315];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[316]; 
@(posedge clk);
#1;data_in = testData6[317];
@(posedge clk);
#1;data_in = testData6[318];
@(posedge clk);
#1;data_in = testData6[319];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[320];
@(posedge clk);
#1;data_in = testData6[321];
@(posedge clk);
#1;data_in = testData6[322];
@(posedge clk);
#1;data_in = testData6[323];
@(posedge clk);
#1;data_in = testData6[324];
@(posedge clk);
#1;data_in = testData6[325];
@(posedge clk);
#1;data_in = testData6[326];
@(posedge clk);
#1;data_in = testData6[327];
@(posedge clk);
#1;data_in = testData6[328];
@(posedge clk);
#1;data_in = testData6[329];
@(posedge clk);
#1;data_in = testData6[330];
@(posedge clk);
#1;data_in = testData6[331];
@(posedge clk);
#1;data_in = testData6[332];
@(posedge clk);
#1;data_in = testData6[333];
@(posedge clk);
#1;data_in = testData6[334];
@(posedge clk);
#1;data_in = testData6[335];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[336]; 
@(posedge clk);
#1;data_in = testData6[337];
@(posedge clk);
#1;data_in = testData6[338];
@(posedge clk);
#1;data_in = testData6[339];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[340];
@(posedge clk);
#1;data_in = testData6[341];
@(posedge clk);
#1;data_in = testData6[342];
@(posedge clk);
#1;data_in = testData6[343];
@(posedge clk);
#1;data_in = testData6[344];
@(posedge clk);
#1;data_in = testData6[345];
@(posedge clk);
#1;data_in = testData6[346];
@(posedge clk);
#1;data_in = testData6[347];
@(posedge clk);
#1;data_in = testData6[348];
@(posedge clk);
#1;data_in = testData6[349];
@(posedge clk);
#1;data_in = testData6[350];
@(posedge clk);
#1;data_in = testData6[351];
@(posedge clk);
#1;data_in = testData6[352];
@(posedge clk);
#1;data_in = testData6[353];
@(posedge clk);
#1;data_in = testData6[354];
@(posedge clk);
#1;data_in = testData6[355];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[356]; 
@(posedge clk);
#1;data_in = testData6[357];
@(posedge clk);
#1;data_in = testData6[358];
@(posedge clk);
#1;data_in = testData6[359];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[360];
@(posedge clk);
#1;data_in = testData6[361];
@(posedge clk);
#1;data_in = testData6[362];
@(posedge clk);
#1;data_in = testData6[363];
@(posedge clk);
#1;data_in = testData6[364];
@(posedge clk);
#1;data_in = testData6[365];
@(posedge clk);
#1;data_in = testData6[366];
@(posedge clk);
#1;data_in = testData6[367];
@(posedge clk);
#1;data_in = testData6[368];
@(posedge clk);
#1;data_in = testData6[369];
@(posedge clk);
#1;data_in = testData6[370];
@(posedge clk);
#1;data_in = testData6[371];
@(posedge clk);
#1;data_in = testData6[372];
@(posedge clk);
#1;data_in = testData6[373];
@(posedge clk);
#1;data_in = testData6[374];
@(posedge clk);
#1;data_in = testData6[375];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[376]; 
@(posedge clk);
#1;data_in = testData6[377];
@(posedge clk);
#1;data_in = testData6[378];
@(posedge clk);
#1;data_in = testData6[379];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[380];
@(posedge clk);
#1;data_in = testData6[381];
@(posedge clk);
#1;data_in = testData6[382];
@(posedge clk);
#1;data_in = testData6[383];
@(posedge clk);
#1;data_in = testData6[384];
@(posedge clk);
#1;data_in = testData6[385];
@(posedge clk);
#1;data_in = testData6[386];
@(posedge clk);
#1;data_in = testData6[387];
@(posedge clk);
#1;data_in = testData6[388];
@(posedge clk);
#1;data_in = testData6[389];
@(posedge clk);
#1;data_in = testData6[390];
@(posedge clk);
#1;data_in = testData6[391];
@(posedge clk);
#1;data_in = testData6[392];
@(posedge clk);
#1;data_in = testData6[393];
@(posedge clk);
#1;data_in = testData6[394];
@(posedge clk);
#1;data_in = testData6[395];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[396]; 
@(posedge clk);
#1;data_in = testData6[397];
@(posedge clk);
#1;data_in = testData6[398];
@(posedge clk);
#1;data_in = testData6[399];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[400];
@(posedge clk);
#1;data_in = testData6[401];
@(posedge clk);
#1;data_in = testData6[402];
@(posedge clk);
#1;data_in = testData6[403];
@(posedge clk);
#1;data_in = testData6[404];
@(posedge clk);
#1;data_in = testData6[405];
@(posedge clk);
#1;data_in = testData6[406];
@(posedge clk);
#1;data_in = testData6[407];
@(posedge clk);
#1;data_in = testData6[408];
@(posedge clk);
#1;data_in = testData6[409];
@(posedge clk);
#1;data_in = testData6[410];
@(posedge clk);
#1;data_in = testData6[411];
@(posedge clk);
#1;data_in = testData6[412];
@(posedge clk);
#1;data_in = testData6[413];
@(posedge clk);
#1;data_in = testData6[414];
@(posedge clk);
#1;data_in = testData6[415];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[416]; 
@(posedge clk);
#1;data_in = testData6[417];
@(posedge clk);
#1;data_in = testData6[418];
@(posedge clk);
#1;data_in = testData6[419];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[420];
@(posedge clk);
#1;data_in = testData6[421];
@(posedge clk);
#1;data_in = testData6[422];
@(posedge clk);
#1;data_in = testData6[423];
@(posedge clk);
#1;data_in = testData6[424];
@(posedge clk);
#1;data_in = testData6[425];
@(posedge clk);
#1;data_in = testData6[426];
@(posedge clk);
#1;data_in = testData6[427];
@(posedge clk);
#1;data_in = testData6[428];
@(posedge clk);
#1;data_in = testData6[429];
@(posedge clk);
#1;data_in = testData6[430];
@(posedge clk);
#1;data_in = testData6[431];
@(posedge clk);
#1;data_in = testData6[432];
@(posedge clk);
#1;data_in = testData6[433];
@(posedge clk);
#1;data_in = testData6[434];
@(posedge clk);
#1;data_in = testData6[435];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[436]; 
@(posedge clk);
#1;data_in = testData6[437];
@(posedge clk);
#1;data_in = testData6[438];
@(posedge clk);
#1;data_in = testData6[439];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[440];
@(posedge clk);
#1;data_in = testData6[441];
@(posedge clk);
#1;data_in = testData6[442];
@(posedge clk);
#1;data_in = testData6[443];
@(posedge clk);
#1;data_in = testData6[444];
@(posedge clk);
#1;data_in = testData6[445];
@(posedge clk);
#1;data_in = testData6[446];
@(posedge clk);
#1;data_in = testData6[447];
@(posedge clk);
#1;data_in = testData6[448];
@(posedge clk);
#1;data_in = testData6[449];
@(posedge clk);
#1;data_in = testData6[450];
@(posedge clk);
#1;data_in = testData6[451];
@(posedge clk);
#1;data_in = testData6[452];
@(posedge clk);
#1;data_in = testData6[453];
@(posedge clk);
#1;data_in = testData6[454];
@(posedge clk);
#1;data_in = testData6[455];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[456]; 
@(posedge clk);
#1;data_in = testData6[457];
@(posedge clk);
#1;data_in = testData6[458];
@(posedge clk);
#1;data_in = testData6[459];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[460];
@(posedge clk);
#1;data_in = testData6[461];
@(posedge clk);
#1;data_in = testData6[462];
@(posedge clk);
#1;data_in = testData6[463];
@(posedge clk);
#1;data_in = testData6[464];
@(posedge clk);
#1;data_in = testData6[465];
@(posedge clk);
#1;data_in = testData6[466];
@(posedge clk);
#1;data_in = testData6[467];
@(posedge clk);
#1;data_in = testData6[468];
@(posedge clk);
#1;data_in = testData6[469];
@(posedge clk);
#1;data_in = testData6[470];
@(posedge clk);
#1;data_in = testData6[471];
@(posedge clk);
#1;data_in = testData6[472];
@(posedge clk);
#1;data_in = testData6[473];
@(posedge clk);
#1;data_in = testData6[474];
@(posedge clk);
#1;data_in = testData6[475];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[476]; 
@(posedge clk);
#1;data_in = testData6[477];
@(posedge clk);
#1;data_in = testData6[478];
@(posedge clk);
#1;data_in = testData6[479];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[480];
@(posedge clk);
#1;data_in = testData6[481];
@(posedge clk);
#1;data_in = testData6[482];
@(posedge clk);
#1;data_in = testData6[483];
@(posedge clk);
#1;data_in = testData6[484];
@(posedge clk);
#1;data_in = testData6[485];
@(posedge clk);
#1;data_in = testData6[486];
@(posedge clk);
#1;data_in = testData6[487];
@(posedge clk);
#1;data_in = testData6[488];
@(posedge clk);
#1;data_in = testData6[489];
@(posedge clk);
#1;data_in = testData6[490];
@(posedge clk);
#1;data_in = testData6[491];
@(posedge clk);
#1;data_in = testData6[492];
@(posedge clk);
#1;data_in = testData6[493];
@(posedge clk);
#1;data_in = testData6[494];
@(posedge clk);
#1;data_in = testData6[495];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[496]; 
@(posedge clk);
#1;data_in = testData6[497];
@(posedge clk);
#1;data_in = testData6[498];
@(posedge clk);
#1;data_in = testData6[499];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[500];
@(posedge clk);
#1;data_in = testData6[501];
@(posedge clk);
#1;data_in = testData6[502];
@(posedge clk);
#1;data_in = testData6[503];
@(posedge clk);
#1;data_in = testData6[504];
@(posedge clk);
#1;data_in = testData6[505];
@(posedge clk);
#1;data_in = testData6[506];
@(posedge clk);
#1;data_in = testData6[507];
@(posedge clk);
#1;data_in = testData6[508];
@(posedge clk);
#1;data_in = testData6[509];
@(posedge clk);
#1;data_in = testData6[510];
@(posedge clk);
#1;data_in = testData6[511];
@(posedge clk);
#1;data_in = testData6[512];
@(posedge clk);
#1;data_in = testData6[513];
@(posedge clk);
#1;data_in = testData6[514];
@(posedge clk);
#1;data_in = testData6[515];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[516]; 
@(posedge clk);
#1;data_in = testData6[517];
@(posedge clk);
#1;data_in = testData6[518];
@(posedge clk);
#1;data_in = testData6[519];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[520];
@(posedge clk);
#1;data_in = testData6[521];
@(posedge clk);
#1;data_in = testData6[522];
@(posedge clk);
#1;data_in = testData6[523];
@(posedge clk);
#1;data_in = testData6[524];
@(posedge clk);
#1;data_in = testData6[525];
@(posedge clk);
#1;data_in = testData6[526];
@(posedge clk);
#1;data_in = testData6[527];
@(posedge clk);
#1;data_in = testData6[528];
@(posedge clk);
#1;data_in = testData6[529];
@(posedge clk);
#1;data_in = testData6[530];
@(posedge clk);
#1;data_in = testData6[531];
@(posedge clk);
#1;data_in = testData6[532];
@(posedge clk);
#1;data_in = testData6[533];
@(posedge clk);
#1;data_in = testData6[534];
@(posedge clk);
#1;data_in = testData6[535];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[536]; 
@(posedge clk);
#1;data_in = testData6[537];
@(posedge clk);
#1;data_in = testData6[538];
@(posedge clk);
#1;data_in = testData6[539];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[540];
@(posedge clk);
#1;data_in = testData6[541];
@(posedge clk);
#1;data_in = testData6[542];
@(posedge clk);
#1;data_in = testData6[543];
@(posedge clk);
#1;data_in = testData6[544];
@(posedge clk);
#1;data_in = testData6[545];
@(posedge clk);
#1;data_in = testData6[546];
@(posedge clk);
#1;data_in = testData6[547];
@(posedge clk);
#1;data_in = testData6[548];
@(posedge clk);
#1;data_in = testData6[549];
@(posedge clk);
#1;data_in = testData6[550];
@(posedge clk);
#1;data_in = testData6[551];
@(posedge clk);
#1;data_in = testData6[552];
@(posedge clk);
#1;data_in = testData6[553];
@(posedge clk);
#1;data_in = testData6[554];
@(posedge clk);
#1;data_in = testData6[555];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[556]; 
@(posedge clk);
#1;data_in = testData6[557];
@(posedge clk);
#1;data_in = testData6[558];
@(posedge clk);
#1;data_in = testData6[559];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[560];
@(posedge clk);
#1;data_in = testData6[561];
@(posedge clk);
#1;data_in = testData6[562];
@(posedge clk);
#1;data_in = testData6[563];
@(posedge clk);
#1;data_in = testData6[564];
@(posedge clk);
#1;data_in = testData6[565];
@(posedge clk);
#1;data_in = testData6[566];
@(posedge clk);
#1;data_in = testData6[567];
@(posedge clk);
#1;data_in = testData6[568];
@(posedge clk);
#1;data_in = testData6[569];
@(posedge clk);
#1;data_in = testData6[570];
@(posedge clk);
#1;data_in = testData6[571];
@(posedge clk);
#1;data_in = testData6[572];
@(posedge clk);
#1;data_in = testData6[573];
@(posedge clk);
#1;data_in = testData6[574];
@(posedge clk);
#1;data_in = testData6[575];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[576]; 
@(posedge clk);
#1;data_in = testData6[577];
@(posedge clk);
#1;data_in = testData6[578];
@(posedge clk);
#1;data_in = testData6[579];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[580];
@(posedge clk);
#1;data_in = testData6[581];
@(posedge clk);
#1;data_in = testData6[582];
@(posedge clk);
#1;data_in = testData6[583];
@(posedge clk);
#1;data_in = testData6[584];
@(posedge clk);
#1;data_in = testData6[585];
@(posedge clk);
#1;data_in = testData6[586];
@(posedge clk);
#1;data_in = testData6[587];
@(posedge clk);
#1;data_in = testData6[588];
@(posedge clk);
#1;data_in = testData6[589];
@(posedge clk);
#1;data_in = testData6[590];
@(posedge clk);
#1;data_in = testData6[591];
@(posedge clk);
#1;data_in = testData6[592];
@(posedge clk);
#1;data_in = testData6[593];
@(posedge clk);
#1;data_in = testData6[594];
@(posedge clk);
#1;data_in = testData6[595];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[596]; 
@(posedge clk);
#1;data_in = testData6[597];
@(posedge clk);
#1;data_in = testData6[598];
@(posedge clk);
#1;data_in = testData6[599];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[600];
@(posedge clk);
#1;data_in = testData6[601];
@(posedge clk);
#1;data_in = testData6[602];
@(posedge clk);
#1;data_in = testData6[603];
@(posedge clk);
#1;data_in = testData6[604];
@(posedge clk);
#1;data_in = testData6[605];
@(posedge clk);
#1;data_in = testData6[606];
@(posedge clk);
#1;data_in = testData6[607];
@(posedge clk);
#1;data_in = testData6[608];
@(posedge clk);
#1;data_in = testData6[609];
@(posedge clk);
#1;data_in = testData6[610];
@(posedge clk);
#1;data_in = testData6[611];
@(posedge clk);
#1;data_in = testData6[612];
@(posedge clk);
#1;data_in = testData6[613];
@(posedge clk);
#1;data_in = testData6[614];
@(posedge clk);
#1;data_in = testData6[615];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[616]; 
@(posedge clk);
#1;data_in = testData6[617];
@(posedge clk);
#1;data_in = testData6[618];
@(posedge clk);
#1;data_in = testData6[619];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[620];
@(posedge clk);
#1;data_in = testData6[621];
@(posedge clk);
#1;data_in = testData6[622];
@(posedge clk);
#1;data_in = testData6[623];
@(posedge clk);
#1;data_in = testData6[624];
@(posedge clk);
#1;data_in = testData6[625];
@(posedge clk);
#1;data_in = testData6[626];
@(posedge clk);
#1;data_in = testData6[627];
@(posedge clk);
#1;data_in = testData6[628];
@(posedge clk);
#1;data_in = testData6[629];
@(posedge clk);
#1;data_in = testData6[630];
@(posedge clk);
#1;data_in = testData6[631];
@(posedge clk);
#1;data_in = testData6[632];
@(posedge clk);
#1;data_in = testData6[633];
@(posedge clk);
#1;data_in = testData6[634];
@(posedge clk);
#1;data_in = testData6[635];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[636]; 
@(posedge clk);
#1;data_in = testData6[637];
@(posedge clk);
#1;data_in = testData6[638];
@(posedge clk);
#1;data_in = testData6[639];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[640];
@(posedge clk);
#1;data_in = testData6[641];
@(posedge clk);
#1;data_in = testData6[642];
@(posedge clk);
#1;data_in = testData6[643];
@(posedge clk);
#1;data_in = testData6[644];
@(posedge clk);
#1;data_in = testData6[645];
@(posedge clk);
#1;data_in = testData6[646];
@(posedge clk);
#1;data_in = testData6[647];
@(posedge clk);
#1;data_in = testData6[648];
@(posedge clk);
#1;data_in = testData6[649];
@(posedge clk);
#1;data_in = testData6[650];
@(posedge clk);
#1;data_in = testData6[651];
@(posedge clk);
#1;data_in = testData6[652];
@(posedge clk);
#1;data_in = testData6[653];
@(posedge clk);
#1;data_in = testData6[654];
@(posedge clk);
#1;data_in = testData6[655];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[656]; 
@(posedge clk);
#1;data_in = testData6[657];
@(posedge clk);
#1;data_in = testData6[658];
@(posedge clk);
#1;data_in = testData6[659];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[660];
@(posedge clk);
#1;data_in = testData6[661];
@(posedge clk);
#1;data_in = testData6[662];
@(posedge clk);
#1;data_in = testData6[663];
@(posedge clk);
#1;data_in = testData6[664];
@(posedge clk);
#1;data_in = testData6[665];
@(posedge clk);
#1;data_in = testData6[666];
@(posedge clk);
#1;data_in = testData6[667];
@(posedge clk);
#1;data_in = testData6[668];
@(posedge clk);
#1;data_in = testData6[669];
@(posedge clk);
#1;data_in = testData6[670];
@(posedge clk);
#1;data_in = testData6[671];
@(posedge clk);
#1;data_in = testData6[672];
@(posedge clk);
#1;data_in = testData6[673];
@(posedge clk);
#1;data_in = testData6[674];
@(posedge clk);
#1;data_in = testData6[675];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[676]; 
@(posedge clk);
#1;data_in = testData6[677];
@(posedge clk);
#1;data_in = testData6[678];
@(posedge clk);
#1;data_in = testData6[679];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[680];
@(posedge clk);
#1;data_in = testData6[681];
@(posedge clk);
#1;data_in = testData6[682];
@(posedge clk);
#1;data_in = testData6[683];
@(posedge clk);
#1;data_in = testData6[684];
@(posedge clk);
#1;data_in = testData6[685];
@(posedge clk);
#1;data_in = testData6[686];
@(posedge clk);
#1;data_in = testData6[687];
@(posedge clk);
#1;data_in = testData6[688];
@(posedge clk);
#1;data_in = testData6[689];
@(posedge clk);
#1;data_in = testData6[690];
@(posedge clk);
#1;data_in = testData6[691];
@(posedge clk);
#1;data_in = testData6[692];
@(posedge clk);
#1;data_in = testData6[693];
@(posedge clk);
#1;data_in = testData6[694];
@(posedge clk);
#1;data_in = testData6[695];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[696]; 
@(posedge clk);
#1;data_in = testData6[697];
@(posedge clk);
#1;data_in = testData6[698];
@(posedge clk);
#1;data_in = testData6[699];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[700];
@(posedge clk);
#1;data_in = testData6[701];
@(posedge clk);
#1;data_in = testData6[702];
@(posedge clk);
#1;data_in = testData6[703];
@(posedge clk);
#1;data_in = testData6[704];
@(posedge clk);
#1;data_in = testData6[705];
@(posedge clk);
#1;data_in = testData6[706];
@(posedge clk);
#1;data_in = testData6[707];
@(posedge clk);
#1;data_in = testData6[708];
@(posedge clk);
#1;data_in = testData6[709];
@(posedge clk);
#1;data_in = testData6[710];
@(posedge clk);
#1;data_in = testData6[711];
@(posedge clk);
#1;data_in = testData6[712];
@(posedge clk);
#1;data_in = testData6[713];
@(posedge clk);
#1;data_in = testData6[714];
@(posedge clk);
#1;data_in = testData6[715];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[716]; 
@(posedge clk);
#1;data_in = testData6[717];
@(posedge clk);
#1;data_in = testData6[718];
@(posedge clk);
#1;data_in = testData6[719];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[720];
@(posedge clk);
#1;data_in = testData6[721];
@(posedge clk);
#1;data_in = testData6[722];
@(posedge clk);
#1;data_in = testData6[723];
@(posedge clk);
#1;data_in = testData6[724];
@(posedge clk);
#1;data_in = testData6[725];
@(posedge clk);
#1;data_in = testData6[726];
@(posedge clk);
#1;data_in = testData6[727];
@(posedge clk);
#1;data_in = testData6[728];
@(posedge clk);
#1;data_in = testData6[729];
@(posedge clk);
#1;data_in = testData6[730];
@(posedge clk);
#1;data_in = testData6[731];
@(posedge clk);
#1;data_in = testData6[732];
@(posedge clk);
#1;data_in = testData6[733];
@(posedge clk);
#1;data_in = testData6[734];
@(posedge clk);
#1;data_in = testData6[735];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[736]; 
@(posedge clk);
#1;data_in = testData6[737];
@(posedge clk);
#1;data_in = testData6[738];
@(posedge clk);
#1;data_in = testData6[739];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[740];
@(posedge clk);
#1;data_in = testData6[741];
@(posedge clk);
#1;data_in = testData6[742];
@(posedge clk);
#1;data_in = testData6[743];
@(posedge clk);
#1;data_in = testData6[744];
@(posedge clk);
#1;data_in = testData6[745];
@(posedge clk);
#1;data_in = testData6[746];
@(posedge clk);
#1;data_in = testData6[747];
@(posedge clk);
#1;data_in = testData6[748];
@(posedge clk);
#1;data_in = testData6[749];
@(posedge clk);
#1;data_in = testData6[750];
@(posedge clk);
#1;data_in = testData6[751];
@(posedge clk);
#1;data_in = testData6[752];
@(posedge clk);
#1;data_in = testData6[753];
@(posedge clk);
#1;data_in = testData6[754];
@(posedge clk);
#1;data_in = testData6[755];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[756]; 
@(posedge clk);
#1;data_in = testData6[757];
@(posedge clk);
#1;data_in = testData6[758];
@(posedge clk);
#1;data_in = testData6[759];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[760];
@(posedge clk);
#1;data_in = testData6[761];
@(posedge clk);
#1;data_in = testData6[762];
@(posedge clk);
#1;data_in = testData6[763];
@(posedge clk);
#1;data_in = testData6[764];
@(posedge clk);
#1;data_in = testData6[765];
@(posedge clk);
#1;data_in = testData6[766];
@(posedge clk);
#1;data_in = testData6[767];
@(posedge clk);
#1;data_in = testData6[768];
@(posedge clk);
#1;data_in = testData6[769];
@(posedge clk);
#1;data_in = testData6[770];
@(posedge clk);
#1;data_in = testData6[771];
@(posedge clk);
#1;data_in = testData6[772];
@(posedge clk);
#1;data_in = testData6[773];
@(posedge clk);
#1;data_in = testData6[774];
@(posedge clk);
#1;data_in = testData6[775];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[776]; 
@(posedge clk);
#1;data_in = testData6[777];
@(posedge clk);
#1;data_in = testData6[778];
@(posedge clk);
#1;data_in = testData6[779];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[780];
@(posedge clk);
#1;data_in = testData6[781];
@(posedge clk);
#1;data_in = testData6[782];
@(posedge clk);
#1;data_in = testData6[783];
@(posedge clk);
#1;data_in = testData6[784];
@(posedge clk);
#1;data_in = testData6[785];
@(posedge clk);
#1;data_in = testData6[786];
@(posedge clk);
#1;data_in = testData6[787];
@(posedge clk);
#1;data_in = testData6[788];
@(posedge clk);
#1;data_in = testData6[789];
@(posedge clk);
#1;data_in = testData6[790];
@(posedge clk);
#1;data_in = testData6[791];
@(posedge clk);
#1;data_in = testData6[792];
@(posedge clk);
#1;data_in = testData6[793];
@(posedge clk);
#1;data_in = testData6[794];
@(posedge clk);
#1;data_in = testData6[795];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[796]; 
@(posedge clk);
#1;data_in = testData6[797];
@(posedge clk);
#1;data_in = testData6[798];
@(posedge clk);
#1;data_in = testData6[799];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[800];
@(posedge clk);
#1;data_in = testData6[801];
@(posedge clk);
#1;data_in = testData6[802];
@(posedge clk);
#1;data_in = testData6[803];
@(posedge clk);
#1;data_in = testData6[804];
@(posedge clk);
#1;data_in = testData6[805];
@(posedge clk);
#1;data_in = testData6[806];
@(posedge clk);
#1;data_in = testData6[807];
@(posedge clk);
#1;data_in = testData6[808];
@(posedge clk);
#1;data_in = testData6[809];
@(posedge clk);
#1;data_in = testData6[810];
@(posedge clk);
#1;data_in = testData6[811];
@(posedge clk);
#1;data_in = testData6[812];
@(posedge clk);
#1;data_in = testData6[813];
@(posedge clk);
#1;data_in = testData6[814];
@(posedge clk);
#1;data_in = testData6[815];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[816]; 
@(posedge clk);
#1;data_in = testData6[817];
@(posedge clk);
#1;data_in = testData6[818];
@(posedge clk);
#1;data_in = testData6[819];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[820];
@(posedge clk);
#1;data_in = testData6[821];
@(posedge clk);
#1;data_in = testData6[822];
@(posedge clk);
#1;data_in = testData6[823];
@(posedge clk);
#1;data_in = testData6[824];
@(posedge clk);
#1;data_in = testData6[825];
@(posedge clk);
#1;data_in = testData6[826];
@(posedge clk);
#1;data_in = testData6[827];
@(posedge clk);
#1;data_in = testData6[828];
@(posedge clk);
#1;data_in = testData6[829];
@(posedge clk);
#1;data_in = testData6[830];
@(posedge clk);
#1;data_in = testData6[831];
@(posedge clk);
#1;data_in = testData6[832];
@(posedge clk);
#1;data_in = testData6[833];
@(posedge clk);
#1;data_in = testData6[834];
@(posedge clk);
#1;data_in = testData6[835];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[836]; 
@(posedge clk);
#1;data_in = testData6[837];
@(posedge clk);
#1;data_in = testData6[838];
@(posedge clk);
#1;data_in = testData6[839];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[840];
@(posedge clk);
#1;data_in = testData6[841];
@(posedge clk);
#1;data_in = testData6[842];
@(posedge clk);
#1;data_in = testData6[843];
@(posedge clk);
#1;data_in = testData6[844];
@(posedge clk);
#1;data_in = testData6[845];
@(posedge clk);
#1;data_in = testData6[846];
@(posedge clk);
#1;data_in = testData6[847];
@(posedge clk);
#1;data_in = testData6[848];
@(posedge clk);
#1;data_in = testData6[849];
@(posedge clk);
#1;data_in = testData6[850];
@(posedge clk);
#1;data_in = testData6[851];
@(posedge clk);
#1;data_in = testData6[852];
@(posedge clk);
#1;data_in = testData6[853];
@(posedge clk);
#1;data_in = testData6[854];
@(posedge clk);
#1;data_in = testData6[855];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[856]; 
@(posedge clk);
#1;data_in = testData6[857];
@(posedge clk);
#1;data_in = testData6[858];
@(posedge clk);
#1;data_in = testData6[859];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[860];
@(posedge clk);
#1;data_in = testData6[861];
@(posedge clk);
#1;data_in = testData6[862];
@(posedge clk);
#1;data_in = testData6[863];
@(posedge clk);
#1;data_in = testData6[864];
@(posedge clk);
#1;data_in = testData6[865];
@(posedge clk);
#1;data_in = testData6[866];
@(posedge clk);
#1;data_in = testData6[867];
@(posedge clk);
#1;data_in = testData6[868];
@(posedge clk);
#1;data_in = testData6[869];
@(posedge clk);
#1;data_in = testData6[870];
@(posedge clk);
#1;data_in = testData6[871];
@(posedge clk);
#1;data_in = testData6[872];
@(posedge clk);
#1;data_in = testData6[873];
@(posedge clk);
#1;data_in = testData6[874];
@(posedge clk);
#1;data_in = testData6[875];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[876]; 
@(posedge clk);
#1;data_in = testData6[877];
@(posedge clk);
#1;data_in = testData6[878];
@(posedge clk);
#1;data_in = testData6[879];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[880];
@(posedge clk);
#1;data_in = testData6[881];
@(posedge clk);
#1;data_in = testData6[882];
@(posedge clk);
#1;data_in = testData6[883];
@(posedge clk);
#1;data_in = testData6[884];
@(posedge clk);
#1;data_in = testData6[885];
@(posedge clk);
#1;data_in = testData6[886];
@(posedge clk);
#1;data_in = testData6[887];
@(posedge clk);
#1;data_in = testData6[888];
@(posedge clk);
#1;data_in = testData6[889];
@(posedge clk);
#1;data_in = testData6[890];
@(posedge clk);
#1;data_in = testData6[891];
@(posedge clk);
#1;data_in = testData6[892];
@(posedge clk);
#1;data_in = testData6[893];
@(posedge clk);
#1;data_in = testData6[894];
@(posedge clk);
#1;data_in = testData6[895];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[896]; 
@(posedge clk);
#1;data_in = testData6[897];
@(posedge clk);
#1;data_in = testData6[898];
@(posedge clk);
#1;data_in = testData6[899];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[900];
@(posedge clk);
#1;data_in = testData6[901];
@(posedge clk);
#1;data_in = testData6[902];
@(posedge clk);
#1;data_in = testData6[903];
@(posedge clk);
#1;data_in = testData6[904];
@(posedge clk);
#1;data_in = testData6[905];
@(posedge clk);
#1;data_in = testData6[906];
@(posedge clk);
#1;data_in = testData6[907];
@(posedge clk);
#1;data_in = testData6[908];
@(posedge clk);
#1;data_in = testData6[909];
@(posedge clk);
#1;data_in = testData6[910];
@(posedge clk);
#1;data_in = testData6[911];
@(posedge clk);
#1;data_in = testData6[912];
@(posedge clk);
#1;data_in = testData6[913];
@(posedge clk);
#1;data_in = testData6[914];
@(posedge clk);
#1;data_in = testData6[915];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[916]; 
@(posedge clk);
#1;data_in = testData6[917];
@(posedge clk);
#1;data_in = testData6[918];
@(posedge clk);
#1;data_in = testData6[919];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[920];
@(posedge clk);
#1;data_in = testData6[921];
@(posedge clk);
#1;data_in = testData6[922];
@(posedge clk);
#1;data_in = testData6[923];
@(posedge clk);
#1;data_in = testData6[924];
@(posedge clk);
#1;data_in = testData6[925];
@(posedge clk);
#1;data_in = testData6[926];
@(posedge clk);
#1;data_in = testData6[927];
@(posedge clk);
#1;data_in = testData6[928];
@(posedge clk);
#1;data_in = testData6[929];
@(posedge clk);
#1;data_in = testData6[930];
@(posedge clk);
#1;data_in = testData6[931];
@(posedge clk);
#1;data_in = testData6[932];
@(posedge clk);
#1;data_in = testData6[933];
@(posedge clk);
#1;data_in = testData6[934];
@(posedge clk);
#1;data_in = testData6[935];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[936]; 
@(posedge clk);
#1;data_in = testData6[937];
@(posedge clk);
#1;data_in = testData6[938];
@(posedge clk);
#1;data_in = testData6[939];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[940];
@(posedge clk);
#1;data_in = testData6[941];
@(posedge clk);
#1;data_in = testData6[942];
@(posedge clk);
#1;data_in = testData6[943];
@(posedge clk);
#1;data_in = testData6[944];
@(posedge clk);
#1;data_in = testData6[945];
@(posedge clk);
#1;data_in = testData6[946];
@(posedge clk);
#1;data_in = testData6[947];
@(posedge clk);
#1;data_in = testData6[948];
@(posedge clk);
#1;data_in = testData6[949];
@(posedge clk);
#1;data_in = testData6[950];
@(posedge clk);
#1;data_in = testData6[951];
@(posedge clk);
#1;data_in = testData6[952];
@(posedge clk);
#1;data_in = testData6[953];
@(posedge clk);
#1;data_in = testData6[954];
@(posedge clk);
#1;data_in = testData6[955];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[956]; 
@(posedge clk);
#1;data_in = testData6[957];
@(posedge clk);
#1;data_in = testData6[958];
@(posedge clk);
#1;data_in = testData6[959];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[960];
@(posedge clk);
#1;data_in = testData6[961];
@(posedge clk);
#1;data_in = testData6[962];
@(posedge clk);
#1;data_in = testData6[963];
@(posedge clk);
#1;data_in = testData6[964];
@(posedge clk);
#1;data_in = testData6[965];
@(posedge clk);
#1;data_in = testData6[966];
@(posedge clk);
#1;data_in = testData6[967];
@(posedge clk);
#1;data_in = testData6[968];
@(posedge clk);
#1;data_in = testData6[969];
@(posedge clk);
#1;data_in = testData6[970];
@(posedge clk);
#1;data_in = testData6[971];
@(posedge clk);
#1;data_in = testData6[972];
@(posedge clk);
#1;data_in = testData6[973];
@(posedge clk);
#1;data_in = testData6[974];
@(posedge clk);
#1;data_in = testData6[975];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[976]; 
@(posedge clk);
#1;data_in = testData6[977];
@(posedge clk);
#1;data_in = testData6[978];
@(posedge clk);
#1;data_in = testData6[979];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[980];
@(posedge clk);
#1;data_in = testData6[981];
@(posedge clk);
#1;data_in = testData6[982];
@(posedge clk);
#1;data_in = testData6[983];
@(posedge clk);
#1;data_in = testData6[984];
@(posedge clk);
#1;data_in = testData6[985];
@(posedge clk);
#1;data_in = testData6[986];
@(posedge clk);
#1;data_in = testData6[987];
@(posedge clk);
#1;data_in = testData6[988];
@(posedge clk);
#1;data_in = testData6[989];
@(posedge clk);
#1;data_in = testData6[990];
@(posedge clk);
#1;data_in = testData6[991];
@(posedge clk);
#1;data_in = testData6[992];
@(posedge clk);
#1;data_in = testData6[993];
@(posedge clk);
#1;data_in = testData6[994];
@(posedge clk);
#1;data_in = testData6[995];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[996]; 
@(posedge clk);
#1;data_in = testData6[997];
@(posedge clk);
#1;data_in = testData6[998];
@(posedge clk);
#1;data_in = testData6[999];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData6[1000];
@(posedge clk);
#1;data_in = testData6[1001];
@(posedge clk);
#1;data_in = testData6[1002];
@(posedge clk);
#1;data_in = testData6[1003];
@(posedge clk);
#1;data_in = testData6[1004];
@(posedge clk);
#1;data_in = testData6[1005];
@(posedge clk);
#1;data_in = testData6[1006];
@(posedge clk);
#1;data_in = testData6[1007];
@(posedge clk);
#1;data_in = testData6[1008];
@(posedge clk);
#1;data_in = testData6[1009];
@(posedge clk);
#1;data_in = testData6[1010];
@(posedge clk);
#1;data_in = testData6[1011];
@(posedge clk);
#1;data_in = testData6[1012];
@(posedge clk);
#1;data_in = testData6[1013];
@(posedge clk);
#1;data_in = testData6[1014];
@(posedge clk);
#1;data_in = testData6[1015];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData6[1016]; 
@(posedge clk);
#1;data_in = testData6[1017];
@(posedge clk);
#1;data_in = testData6[1018];
@(posedge clk);
#1;data_in = testData6[1019];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;

// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
// Testbench, with parameters k=4, p=4, b=8, g=1

module tb5();
logic clk, reset, start, done,qwerty, loadMatrix, loadVector;
 
logic signed [7:0] data_in;
logic signed [15:0] data_out;
mvm_4_4_8_1 dut(clk, reset, loadMatrix, loadVector, start, done, data_in, data_out);

initial clk=0;
   always #5 clk = ~clk;;

logic [7:0] testData5[819:0];
   //read input from C file inputDatapart1     
 initial $readmemh("proj3_inputDatatb5", testData5);
 integer i;
 integer filehandle=$fopen("proj3_outValuestb5");
  initial begin 
  $monitor("Data in : %x",data_in);       
start  = 0; reset  = 1; data_in = 8'bx;
 @(posedge clk); #1; reset=0; loadMatrix=1;      
@(posedge clk);
#1; loadMatrix=0; data_in = testData5[0];
@(posedge clk);
#1;data_in = testData5[1];
@(posedge clk);
#1;data_in = testData5[2];
@(posedge clk);
#1;data_in = testData5[3];
@(posedge clk);
#1;data_in = testData5[4];
@(posedge clk);
#1;data_in = testData5[5];
@(posedge clk);
#1;data_in = testData5[6];
@(posedge clk);
#1;data_in = testData5[7];
@(posedge clk);
#1;data_in = testData5[8];
@(posedge clk);
#1;data_in = testData5[9];
@(posedge clk);
#1;data_in = testData5[10];
@(posedge clk);
#1;data_in = testData5[11];
@(posedge clk);
#1;data_in = testData5[12];
@(posedge clk);
#1;data_in = testData5[13];
@(posedge clk);
#1;data_in = testData5[14];
@(posedge clk);
#1;data_in = testData5[15];
@(posedge clk);
#1; loadVector=1; 
@(posedge clk);
#1; loadVector=0; data_in=testData5[16]; 
@(posedge clk);
#1;data_in = testData5[17];
@(posedge clk);
#1;data_in = testData5[18];
@(posedge clk);
#1;data_in = testData5[19];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[20]; 
@(posedge clk);
#1;data_in = testData5[21];
@(posedge clk);
#1;data_in = testData5[22];
@(posedge clk);
#1;data_in = testData5[23];
@(posedge clk);
#1;data_in = testData5[24];
@(posedge clk);
#1;data_in = testData5[25];
@(posedge clk);
#1;data_in = testData5[26];
@(posedge clk);
#1;data_in = testData5[27];
@(posedge clk);
#1;data_in = testData5[28];
@(posedge clk);
#1;data_in = testData5[29];
@(posedge clk);
#1;data_in = testData5[30];
@(posedge clk);
#1;data_in = testData5[31];
@(posedge clk);
#1;data_in = testData5[32];
@(posedge clk);
#1;data_in = testData5[33];
@(posedge clk);
#1;data_in = testData5[34];
@(posedge clk);
#1;data_in = testData5[35];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[36]; 
@(posedge clk);
#1;data_in = testData5[37];
@(posedge clk);
#1;data_in = testData5[38];
@(posedge clk);
#1;data_in = testData5[39];
@(posedge clk);
#1;data_in = testData5[40];
@(posedge clk);
#1;data_in = testData5[41];
@(posedge clk);
#1;data_in = testData5[42];
@(posedge clk);
#1;data_in = testData5[43];
@(posedge clk);
#1;data_in = testData5[44];
@(posedge clk);
#1;data_in = testData5[45];
@(posedge clk);
#1;data_in = testData5[46];
@(posedge clk);
#1;data_in = testData5[47];
@(posedge clk);
#1;data_in = testData5[48];
@(posedge clk);
#1;data_in = testData5[49];
@(posedge clk);
#1;data_in = testData5[50];
@(posedge clk);
#1;data_in = testData5[51];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[52]; 
@(posedge clk);
#1;data_in = testData5[53];
@(posedge clk);
#1;data_in = testData5[54];
@(posedge clk);
#1;data_in = testData5[55];
@(posedge clk);
#1;data_in = testData5[56];
@(posedge clk);
#1;data_in = testData5[57];
@(posedge clk);
#1;data_in = testData5[58];
@(posedge clk);
#1;data_in = testData5[59];
@(posedge clk);
#1;data_in = testData5[60];
@(posedge clk);
#1;data_in = testData5[61];
@(posedge clk);
#1;data_in = testData5[62];
@(posedge clk);
#1;data_in = testData5[63];
@(posedge clk);
#1;data_in = testData5[64];
@(posedge clk);
#1;data_in = testData5[65];
@(posedge clk);
#1;data_in = testData5[66];
@(posedge clk);
#1;data_in = testData5[67];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[68]; 
@(posedge clk);
#1;data_in = testData5[69];
@(posedge clk);
#1;data_in = testData5[70];
@(posedge clk);
#1;data_in = testData5[71];
@(posedge clk);
#1;data_in = testData5[72];
@(posedge clk);
#1;data_in = testData5[73];
@(posedge clk);
#1;data_in = testData5[74];
@(posedge clk);
#1;data_in = testData5[75];
@(posedge clk);
#1;data_in = testData5[76];
@(posedge clk);
#1;data_in = testData5[77];
@(posedge clk);
#1;data_in = testData5[78];
@(posedge clk);
#1;data_in = testData5[79];
@(posedge clk);
#1;data_in = testData5[80];
@(posedge clk);
#1;data_in = testData5[81];
@(posedge clk);
#1;data_in = testData5[82];
@(posedge clk);
#1;data_in = testData5[83];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[84]; 
@(posedge clk);
#1;data_in = testData5[85];
@(posedge clk);
#1;data_in = testData5[86];
@(posedge clk);
#1;data_in = testData5[87];
@(posedge clk);
#1;data_in = testData5[88];
@(posedge clk);
#1;data_in = testData5[89];
@(posedge clk);
#1;data_in = testData5[90];
@(posedge clk);
#1;data_in = testData5[91];
@(posedge clk);
#1;data_in = testData5[92];
@(posedge clk);
#1;data_in = testData5[93];
@(posedge clk);
#1;data_in = testData5[94];
@(posedge clk);
#1;data_in = testData5[95];
@(posedge clk);
#1;data_in = testData5[96];
@(posedge clk);
#1;data_in = testData5[97];
@(posedge clk);
#1;data_in = testData5[98];
@(posedge clk);
#1;data_in = testData5[99];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[100]; 
@(posedge clk);
#1;data_in = testData5[101];
@(posedge clk);
#1;data_in = testData5[102];
@(posedge clk);
#1;data_in = testData5[103];
@(posedge clk);
#1;data_in = testData5[104];
@(posedge clk);
#1;data_in = testData5[105];
@(posedge clk);
#1;data_in = testData5[106];
@(posedge clk);
#1;data_in = testData5[107];
@(posedge clk);
#1;data_in = testData5[108];
@(posedge clk);
#1;data_in = testData5[109];
@(posedge clk);
#1;data_in = testData5[110];
@(posedge clk);
#1;data_in = testData5[111];
@(posedge clk);
#1;data_in = testData5[112];
@(posedge clk);
#1;data_in = testData5[113];
@(posedge clk);
#1;data_in = testData5[114];
@(posedge clk);
#1;data_in = testData5[115];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[116]; 
@(posedge clk);
#1;data_in = testData5[117];
@(posedge clk);
#1;data_in = testData5[118];
@(posedge clk);
#1;data_in = testData5[119];
@(posedge clk);
#1;data_in = testData5[120];
@(posedge clk);
#1;data_in = testData5[121];
@(posedge clk);
#1;data_in = testData5[122];
@(posedge clk);
#1;data_in = testData5[123];
@(posedge clk);
#1;data_in = testData5[124];
@(posedge clk);
#1;data_in = testData5[125];
@(posedge clk);
#1;data_in = testData5[126];
@(posedge clk);
#1;data_in = testData5[127];
@(posedge clk);
#1;data_in = testData5[128];
@(posedge clk);
#1;data_in = testData5[129];
@(posedge clk);
#1;data_in = testData5[130];
@(posedge clk);
#1;data_in = testData5[131];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[132]; 
@(posedge clk);
#1;data_in = testData5[133];
@(posedge clk);
#1;data_in = testData5[134];
@(posedge clk);
#1;data_in = testData5[135];
@(posedge clk);
#1;data_in = testData5[136];
@(posedge clk);
#1;data_in = testData5[137];
@(posedge clk);
#1;data_in = testData5[138];
@(posedge clk);
#1;data_in = testData5[139];
@(posedge clk);
#1;data_in = testData5[140];
@(posedge clk);
#1;data_in = testData5[141];
@(posedge clk);
#1;data_in = testData5[142];
@(posedge clk);
#1;data_in = testData5[143];
@(posedge clk);
#1;data_in = testData5[144];
@(posedge clk);
#1;data_in = testData5[145];
@(posedge clk);
#1;data_in = testData5[146];
@(posedge clk);
#1;data_in = testData5[147];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[148]; 
@(posedge clk);
#1;data_in = testData5[149];
@(posedge clk);
#1;data_in = testData5[150];
@(posedge clk);
#1;data_in = testData5[151];
@(posedge clk);
#1;data_in = testData5[152];
@(posedge clk);
#1;data_in = testData5[153];
@(posedge clk);
#1;data_in = testData5[154];
@(posedge clk);
#1;data_in = testData5[155];
@(posedge clk);
#1;data_in = testData5[156];
@(posedge clk);
#1;data_in = testData5[157];
@(posedge clk);
#1;data_in = testData5[158];
@(posedge clk);
#1;data_in = testData5[159];
@(posedge clk);
#1;data_in = testData5[160];
@(posedge clk);
#1;data_in = testData5[161];
@(posedge clk);
#1;data_in = testData5[162];
@(posedge clk);
#1;data_in = testData5[163];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[164]; 
@(posedge clk);
#1;data_in = testData5[165];
@(posedge clk);
#1;data_in = testData5[166];
@(posedge clk);
#1;data_in = testData5[167];
@(posedge clk);
#1;data_in = testData5[168];
@(posedge clk);
#1;data_in = testData5[169];
@(posedge clk);
#1;data_in = testData5[170];
@(posedge clk);
#1;data_in = testData5[171];
@(posedge clk);
#1;data_in = testData5[172];
@(posedge clk);
#1;data_in = testData5[173];
@(posedge clk);
#1;data_in = testData5[174];
@(posedge clk);
#1;data_in = testData5[175];
@(posedge clk);
#1;data_in = testData5[176];
@(posedge clk);
#1;data_in = testData5[177];
@(posedge clk);
#1;data_in = testData5[178];
@(posedge clk);
#1;data_in = testData5[179];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[180]; 
@(posedge clk);
#1;data_in = testData5[181];
@(posedge clk);
#1;data_in = testData5[182];
@(posedge clk);
#1;data_in = testData5[183];
@(posedge clk);
#1;data_in = testData5[184];
@(posedge clk);
#1;data_in = testData5[185];
@(posedge clk);
#1;data_in = testData5[186];
@(posedge clk);
#1;data_in = testData5[187];
@(posedge clk);
#1;data_in = testData5[188];
@(posedge clk);
#1;data_in = testData5[189];
@(posedge clk);
#1;data_in = testData5[190];
@(posedge clk);
#1;data_in = testData5[191];
@(posedge clk);
#1;data_in = testData5[192];
@(posedge clk);
#1;data_in = testData5[193];
@(posedge clk);
#1;data_in = testData5[194];
@(posedge clk);
#1;data_in = testData5[195];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[196]; 
@(posedge clk);
#1;data_in = testData5[197];
@(posedge clk);
#1;data_in = testData5[198];
@(posedge clk);
#1;data_in = testData5[199];
@(posedge clk);
#1;data_in = testData5[200];
@(posedge clk);
#1;data_in = testData5[201];
@(posedge clk);
#1;data_in = testData5[202];
@(posedge clk);
#1;data_in = testData5[203];
@(posedge clk);
#1;data_in = testData5[204];
@(posedge clk);
#1;data_in = testData5[205];
@(posedge clk);
#1;data_in = testData5[206];
@(posedge clk);
#1;data_in = testData5[207];
@(posedge clk);
#1;data_in = testData5[208];
@(posedge clk);
#1;data_in = testData5[209];
@(posedge clk);
#1;data_in = testData5[210];
@(posedge clk);
#1;data_in = testData5[211];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[212]; 
@(posedge clk);
#1;data_in = testData5[213];
@(posedge clk);
#1;data_in = testData5[214];
@(posedge clk);
#1;data_in = testData5[215];
@(posedge clk);
#1;data_in = testData5[216];
@(posedge clk);
#1;data_in = testData5[217];
@(posedge clk);
#1;data_in = testData5[218];
@(posedge clk);
#1;data_in = testData5[219];
@(posedge clk);
#1;data_in = testData5[220];
@(posedge clk);
#1;data_in = testData5[221];
@(posedge clk);
#1;data_in = testData5[222];
@(posedge clk);
#1;data_in = testData5[223];
@(posedge clk);
#1;data_in = testData5[224];
@(posedge clk);
#1;data_in = testData5[225];
@(posedge clk);
#1;data_in = testData5[226];
@(posedge clk);
#1;data_in = testData5[227];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[228]; 
@(posedge clk);
#1;data_in = testData5[229];
@(posedge clk);
#1;data_in = testData5[230];
@(posedge clk);
#1;data_in = testData5[231];
@(posedge clk);
#1;data_in = testData5[232];
@(posedge clk);
#1;data_in = testData5[233];
@(posedge clk);
#1;data_in = testData5[234];
@(posedge clk);
#1;data_in = testData5[235];
@(posedge clk);
#1;data_in = testData5[236];
@(posedge clk);
#1;data_in = testData5[237];
@(posedge clk);
#1;data_in = testData5[238];
@(posedge clk);
#1;data_in = testData5[239];
@(posedge clk);
#1;data_in = testData5[240];
@(posedge clk);
#1;data_in = testData5[241];
@(posedge clk);
#1;data_in = testData5[242];
@(posedge clk);
#1;data_in = testData5[243];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[244]; 
@(posedge clk);
#1;data_in = testData5[245];
@(posedge clk);
#1;data_in = testData5[246];
@(posedge clk);
#1;data_in = testData5[247];
@(posedge clk);
#1;data_in = testData5[248];
@(posedge clk);
#1;data_in = testData5[249];
@(posedge clk);
#1;data_in = testData5[250];
@(posedge clk);
#1;data_in = testData5[251];
@(posedge clk);
#1;data_in = testData5[252];
@(posedge clk);
#1;data_in = testData5[253];
@(posedge clk);
#1;data_in = testData5[254];
@(posedge clk);
#1;data_in = testData5[255];
@(posedge clk);
#1;data_in = testData5[256];
@(posedge clk);
#1;data_in = testData5[257];
@(posedge clk);
#1;data_in = testData5[258];
@(posedge clk);
#1;data_in = testData5[259];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[260]; 
@(posedge clk);
#1;data_in = testData5[261];
@(posedge clk);
#1;data_in = testData5[262];
@(posedge clk);
#1;data_in = testData5[263];
@(posedge clk);
#1;data_in = testData5[264];
@(posedge clk);
#1;data_in = testData5[265];
@(posedge clk);
#1;data_in = testData5[266];
@(posedge clk);
#1;data_in = testData5[267];
@(posedge clk);
#1;data_in = testData5[268];
@(posedge clk);
#1;data_in = testData5[269];
@(posedge clk);
#1;data_in = testData5[270];
@(posedge clk);
#1;data_in = testData5[271];
@(posedge clk);
#1;data_in = testData5[272];
@(posedge clk);
#1;data_in = testData5[273];
@(posedge clk);
#1;data_in = testData5[274];
@(posedge clk);
#1;data_in = testData5[275];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[276]; 
@(posedge clk);
#1;data_in = testData5[277];
@(posedge clk);
#1;data_in = testData5[278];
@(posedge clk);
#1;data_in = testData5[279];
@(posedge clk);
#1;data_in = testData5[280];
@(posedge clk);
#1;data_in = testData5[281];
@(posedge clk);
#1;data_in = testData5[282];
@(posedge clk);
#1;data_in = testData5[283];
@(posedge clk);
#1;data_in = testData5[284];
@(posedge clk);
#1;data_in = testData5[285];
@(posedge clk);
#1;data_in = testData5[286];
@(posedge clk);
#1;data_in = testData5[287];
@(posedge clk);
#1;data_in = testData5[288];
@(posedge clk);
#1;data_in = testData5[289];
@(posedge clk);
#1;data_in = testData5[290];
@(posedge clk);
#1;data_in = testData5[291];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[292]; 
@(posedge clk);
#1;data_in = testData5[293];
@(posedge clk);
#1;data_in = testData5[294];
@(posedge clk);
#1;data_in = testData5[295];
@(posedge clk);
#1;data_in = testData5[296];
@(posedge clk);
#1;data_in = testData5[297];
@(posedge clk);
#1;data_in = testData5[298];
@(posedge clk);
#1;data_in = testData5[299];
@(posedge clk);
#1;data_in = testData5[300];
@(posedge clk);
#1;data_in = testData5[301];
@(posedge clk);
#1;data_in = testData5[302];
@(posedge clk);
#1;data_in = testData5[303];
@(posedge clk);
#1;data_in = testData5[304];
@(posedge clk);
#1;data_in = testData5[305];
@(posedge clk);
#1;data_in = testData5[306];
@(posedge clk);
#1;data_in = testData5[307];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[308]; 
@(posedge clk);
#1;data_in = testData5[309];
@(posedge clk);
#1;data_in = testData5[310];
@(posedge clk);
#1;data_in = testData5[311];
@(posedge clk);
#1;data_in = testData5[312];
@(posedge clk);
#1;data_in = testData5[313];
@(posedge clk);
#1;data_in = testData5[314];
@(posedge clk);
#1;data_in = testData5[315];
@(posedge clk);
#1;data_in = testData5[316];
@(posedge clk);
#1;data_in = testData5[317];
@(posedge clk);
#1;data_in = testData5[318];
@(posedge clk);
#1;data_in = testData5[319];
@(posedge clk);
#1;data_in = testData5[320];
@(posedge clk);
#1;data_in = testData5[321];
@(posedge clk);
#1;data_in = testData5[322];
@(posedge clk);
#1;data_in = testData5[323];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[324]; 
@(posedge clk);
#1;data_in = testData5[325];
@(posedge clk);
#1;data_in = testData5[326];
@(posedge clk);
#1;data_in = testData5[327];
@(posedge clk);
#1;data_in = testData5[328];
@(posedge clk);
#1;data_in = testData5[329];
@(posedge clk);
#1;data_in = testData5[330];
@(posedge clk);
#1;data_in = testData5[331];
@(posedge clk);
#1;data_in = testData5[332];
@(posedge clk);
#1;data_in = testData5[333];
@(posedge clk);
#1;data_in = testData5[334];
@(posedge clk);
#1;data_in = testData5[335];
@(posedge clk);
#1;data_in = testData5[336];
@(posedge clk);
#1;data_in = testData5[337];
@(posedge clk);
#1;data_in = testData5[338];
@(posedge clk);
#1;data_in = testData5[339];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[340]; 
@(posedge clk);
#1;data_in = testData5[341];
@(posedge clk);
#1;data_in = testData5[342];
@(posedge clk);
#1;data_in = testData5[343];
@(posedge clk);
#1;data_in = testData5[344];
@(posedge clk);
#1;data_in = testData5[345];
@(posedge clk);
#1;data_in = testData5[346];
@(posedge clk);
#1;data_in = testData5[347];
@(posedge clk);
#1;data_in = testData5[348];
@(posedge clk);
#1;data_in = testData5[349];
@(posedge clk);
#1;data_in = testData5[350];
@(posedge clk);
#1;data_in = testData5[351];
@(posedge clk);
#1;data_in = testData5[352];
@(posedge clk);
#1;data_in = testData5[353];
@(posedge clk);
#1;data_in = testData5[354];
@(posedge clk);
#1;data_in = testData5[355];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[356]; 
@(posedge clk);
#1;data_in = testData5[357];
@(posedge clk);
#1;data_in = testData5[358];
@(posedge clk);
#1;data_in = testData5[359];
@(posedge clk);
#1;data_in = testData5[360];
@(posedge clk);
#1;data_in = testData5[361];
@(posedge clk);
#1;data_in = testData5[362];
@(posedge clk);
#1;data_in = testData5[363];
@(posedge clk);
#1;data_in = testData5[364];
@(posedge clk);
#1;data_in = testData5[365];
@(posedge clk);
#1;data_in = testData5[366];
@(posedge clk);
#1;data_in = testData5[367];
@(posedge clk);
#1;data_in = testData5[368];
@(posedge clk);
#1;data_in = testData5[369];
@(posedge clk);
#1;data_in = testData5[370];
@(posedge clk);
#1;data_in = testData5[371];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[372]; 
@(posedge clk);
#1;data_in = testData5[373];
@(posedge clk);
#1;data_in = testData5[374];
@(posedge clk);
#1;data_in = testData5[375];
@(posedge clk);
#1;data_in = testData5[376];
@(posedge clk);
#1;data_in = testData5[377];
@(posedge clk);
#1;data_in = testData5[378];
@(posedge clk);
#1;data_in = testData5[379];
@(posedge clk);
#1;data_in = testData5[380];
@(posedge clk);
#1;data_in = testData5[381];
@(posedge clk);
#1;data_in = testData5[382];
@(posedge clk);
#1;data_in = testData5[383];
@(posedge clk);
#1;data_in = testData5[384];
@(posedge clk);
#1;data_in = testData5[385];
@(posedge clk);
#1;data_in = testData5[386];
@(posedge clk);
#1;data_in = testData5[387];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[388]; 
@(posedge clk);
#1;data_in = testData5[389];
@(posedge clk);
#1;data_in = testData5[390];
@(posedge clk);
#1;data_in = testData5[391];
@(posedge clk);
#1;data_in = testData5[392];
@(posedge clk);
#1;data_in = testData5[393];
@(posedge clk);
#1;data_in = testData5[394];
@(posedge clk);
#1;data_in = testData5[395];
@(posedge clk);
#1;data_in = testData5[396];
@(posedge clk);
#1;data_in = testData5[397];
@(posedge clk);
#1;data_in = testData5[398];
@(posedge clk);
#1;data_in = testData5[399];
@(posedge clk);
#1;data_in = testData5[400];
@(posedge clk);
#1;data_in = testData5[401];
@(posedge clk);
#1;data_in = testData5[402];
@(posedge clk);
#1;data_in = testData5[403];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[404]; 
@(posedge clk);
#1;data_in = testData5[405];
@(posedge clk);
#1;data_in = testData5[406];
@(posedge clk);
#1;data_in = testData5[407];
@(posedge clk);
#1;data_in = testData5[408];
@(posedge clk);
#1;data_in = testData5[409];
@(posedge clk);
#1;data_in = testData5[410];
@(posedge clk);
#1;data_in = testData5[411];
@(posedge clk);
#1;data_in = testData5[412];
@(posedge clk);
#1;data_in = testData5[413];
@(posedge clk);
#1;data_in = testData5[414];
@(posedge clk);
#1;data_in = testData5[415];
@(posedge clk);
#1;data_in = testData5[416];
@(posedge clk);
#1;data_in = testData5[417];
@(posedge clk);
#1;data_in = testData5[418];
@(posedge clk);
#1;data_in = testData5[419];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[420]; 
@(posedge clk);
#1;data_in = testData5[421];
@(posedge clk);
#1;data_in = testData5[422];
@(posedge clk);
#1;data_in = testData5[423];
@(posedge clk);
#1;data_in = testData5[424];
@(posedge clk);
#1;data_in = testData5[425];
@(posedge clk);
#1;data_in = testData5[426];
@(posedge clk);
#1;data_in = testData5[427];
@(posedge clk);
#1;data_in = testData5[428];
@(posedge clk);
#1;data_in = testData5[429];
@(posedge clk);
#1;data_in = testData5[430];
@(posedge clk);
#1;data_in = testData5[431];
@(posedge clk);
#1;data_in = testData5[432];
@(posedge clk);
#1;data_in = testData5[433];
@(posedge clk);
#1;data_in = testData5[434];
@(posedge clk);
#1;data_in = testData5[435];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[436]; 
@(posedge clk);
#1;data_in = testData5[437];
@(posedge clk);
#1;data_in = testData5[438];
@(posedge clk);
#1;data_in = testData5[439];
@(posedge clk);
#1;data_in = testData5[440];
@(posedge clk);
#1;data_in = testData5[441];
@(posedge clk);
#1;data_in = testData5[442];
@(posedge clk);
#1;data_in = testData5[443];
@(posedge clk);
#1;data_in = testData5[444];
@(posedge clk);
#1;data_in = testData5[445];
@(posedge clk);
#1;data_in = testData5[446];
@(posedge clk);
#1;data_in = testData5[447];
@(posedge clk);
#1;data_in = testData5[448];
@(posedge clk);
#1;data_in = testData5[449];
@(posedge clk);
#1;data_in = testData5[450];
@(posedge clk);
#1;data_in = testData5[451];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[452]; 
@(posedge clk);
#1;data_in = testData5[453];
@(posedge clk);
#1;data_in = testData5[454];
@(posedge clk);
#1;data_in = testData5[455];
@(posedge clk);
#1;data_in = testData5[456];
@(posedge clk);
#1;data_in = testData5[457];
@(posedge clk);
#1;data_in = testData5[458];
@(posedge clk);
#1;data_in = testData5[459];
@(posedge clk);
#1;data_in = testData5[460];
@(posedge clk);
#1;data_in = testData5[461];
@(posedge clk);
#1;data_in = testData5[462];
@(posedge clk);
#1;data_in = testData5[463];
@(posedge clk);
#1;data_in = testData5[464];
@(posedge clk);
#1;data_in = testData5[465];
@(posedge clk);
#1;data_in = testData5[466];
@(posedge clk);
#1;data_in = testData5[467];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[468]; 
@(posedge clk);
#1;data_in = testData5[469];
@(posedge clk);
#1;data_in = testData5[470];
@(posedge clk);
#1;data_in = testData5[471];
@(posedge clk);
#1;data_in = testData5[472];
@(posedge clk);
#1;data_in = testData5[473];
@(posedge clk);
#1;data_in = testData5[474];
@(posedge clk);
#1;data_in = testData5[475];
@(posedge clk);
#1;data_in = testData5[476];
@(posedge clk);
#1;data_in = testData5[477];
@(posedge clk);
#1;data_in = testData5[478];
@(posedge clk);
#1;data_in = testData5[479];
@(posedge clk);
#1;data_in = testData5[480];
@(posedge clk);
#1;data_in = testData5[481];
@(posedge clk);
#1;data_in = testData5[482];
@(posedge clk);
#1;data_in = testData5[483];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[484]; 
@(posedge clk);
#1;data_in = testData5[485];
@(posedge clk);
#1;data_in = testData5[486];
@(posedge clk);
#1;data_in = testData5[487];
@(posedge clk);
#1;data_in = testData5[488];
@(posedge clk);
#1;data_in = testData5[489];
@(posedge clk);
#1;data_in = testData5[490];
@(posedge clk);
#1;data_in = testData5[491];
@(posedge clk);
#1;data_in = testData5[492];
@(posedge clk);
#1;data_in = testData5[493];
@(posedge clk);
#1;data_in = testData5[494];
@(posedge clk);
#1;data_in = testData5[495];
@(posedge clk);
#1;data_in = testData5[496];
@(posedge clk);
#1;data_in = testData5[497];
@(posedge clk);
#1;data_in = testData5[498];
@(posedge clk);
#1;data_in = testData5[499];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[500]; 
@(posedge clk);
#1;data_in = testData5[501];
@(posedge clk);
#1;data_in = testData5[502];
@(posedge clk);
#1;data_in = testData5[503];
@(posedge clk);
#1;data_in = testData5[504];
@(posedge clk);
#1;data_in = testData5[505];
@(posedge clk);
#1;data_in = testData5[506];
@(posedge clk);
#1;data_in = testData5[507];
@(posedge clk);
#1;data_in = testData5[508];
@(posedge clk);
#1;data_in = testData5[509];
@(posedge clk);
#1;data_in = testData5[510];
@(posedge clk);
#1;data_in = testData5[511];
@(posedge clk);
#1;data_in = testData5[512];
@(posedge clk);
#1;data_in = testData5[513];
@(posedge clk);
#1;data_in = testData5[514];
@(posedge clk);
#1;data_in = testData5[515];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[516]; 
@(posedge clk);
#1;data_in = testData5[517];
@(posedge clk);
#1;data_in = testData5[518];
@(posedge clk);
#1;data_in = testData5[519];
@(posedge clk);
#1;data_in = testData5[520];
@(posedge clk);
#1;data_in = testData5[521];
@(posedge clk);
#1;data_in = testData5[522];
@(posedge clk);
#1;data_in = testData5[523];
@(posedge clk);
#1;data_in = testData5[524];
@(posedge clk);
#1;data_in = testData5[525];
@(posedge clk);
#1;data_in = testData5[526];
@(posedge clk);
#1;data_in = testData5[527];
@(posedge clk);
#1;data_in = testData5[528];
@(posedge clk);
#1;data_in = testData5[529];
@(posedge clk);
#1;data_in = testData5[530];
@(posedge clk);
#1;data_in = testData5[531];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[532]; 
@(posedge clk);
#1;data_in = testData5[533];
@(posedge clk);
#1;data_in = testData5[534];
@(posedge clk);
#1;data_in = testData5[535];
@(posedge clk);
#1;data_in = testData5[536];
@(posedge clk);
#1;data_in = testData5[537];
@(posedge clk);
#1;data_in = testData5[538];
@(posedge clk);
#1;data_in = testData5[539];
@(posedge clk);
#1;data_in = testData5[540];
@(posedge clk);
#1;data_in = testData5[541];
@(posedge clk);
#1;data_in = testData5[542];
@(posedge clk);
#1;data_in = testData5[543];
@(posedge clk);
#1;data_in = testData5[544];
@(posedge clk);
#1;data_in = testData5[545];
@(posedge clk);
#1;data_in = testData5[546];
@(posedge clk);
#1;data_in = testData5[547];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[548]; 
@(posedge clk);
#1;data_in = testData5[549];
@(posedge clk);
#1;data_in = testData5[550];
@(posedge clk);
#1;data_in = testData5[551];
@(posedge clk);
#1;data_in = testData5[552];
@(posedge clk);
#1;data_in = testData5[553];
@(posedge clk);
#1;data_in = testData5[554];
@(posedge clk);
#1;data_in = testData5[555];
@(posedge clk);
#1;data_in = testData5[556];
@(posedge clk);
#1;data_in = testData5[557];
@(posedge clk);
#1;data_in = testData5[558];
@(posedge clk);
#1;data_in = testData5[559];
@(posedge clk);
#1;data_in = testData5[560];
@(posedge clk);
#1;data_in = testData5[561];
@(posedge clk);
#1;data_in = testData5[562];
@(posedge clk);
#1;data_in = testData5[563];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[564]; 
@(posedge clk);
#1;data_in = testData5[565];
@(posedge clk);
#1;data_in = testData5[566];
@(posedge clk);
#1;data_in = testData5[567];
@(posedge clk);
#1;data_in = testData5[568];
@(posedge clk);
#1;data_in = testData5[569];
@(posedge clk);
#1;data_in = testData5[570];
@(posedge clk);
#1;data_in = testData5[571];
@(posedge clk);
#1;data_in = testData5[572];
@(posedge clk);
#1;data_in = testData5[573];
@(posedge clk);
#1;data_in = testData5[574];
@(posedge clk);
#1;data_in = testData5[575];
@(posedge clk);
#1;data_in = testData5[576];
@(posedge clk);
#1;data_in = testData5[577];
@(posedge clk);
#1;data_in = testData5[578];
@(posedge clk);
#1;data_in = testData5[579];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[580]; 
@(posedge clk);
#1;data_in = testData5[581];
@(posedge clk);
#1;data_in = testData5[582];
@(posedge clk);
#1;data_in = testData5[583];
@(posedge clk);
#1;data_in = testData5[584];
@(posedge clk);
#1;data_in = testData5[585];
@(posedge clk);
#1;data_in = testData5[586];
@(posedge clk);
#1;data_in = testData5[587];
@(posedge clk);
#1;data_in = testData5[588];
@(posedge clk);
#1;data_in = testData5[589];
@(posedge clk);
#1;data_in = testData5[590];
@(posedge clk);
#1;data_in = testData5[591];
@(posedge clk);
#1;data_in = testData5[592];
@(posedge clk);
#1;data_in = testData5[593];
@(posedge clk);
#1;data_in = testData5[594];
@(posedge clk);
#1;data_in = testData5[595];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[596]; 
@(posedge clk);
#1;data_in = testData5[597];
@(posedge clk);
#1;data_in = testData5[598];
@(posedge clk);
#1;data_in = testData5[599];
@(posedge clk);
#1;data_in = testData5[600];
@(posedge clk);
#1;data_in = testData5[601];
@(posedge clk);
#1;data_in = testData5[602];
@(posedge clk);
#1;data_in = testData5[603];
@(posedge clk);
#1;data_in = testData5[604];
@(posedge clk);
#1;data_in = testData5[605];
@(posedge clk);
#1;data_in = testData5[606];
@(posedge clk);
#1;data_in = testData5[607];
@(posedge clk);
#1;data_in = testData5[608];
@(posedge clk);
#1;data_in = testData5[609];
@(posedge clk);
#1;data_in = testData5[610];
@(posedge clk);
#1;data_in = testData5[611];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[612]; 
@(posedge clk);
#1;data_in = testData5[613];
@(posedge clk);
#1;data_in = testData5[614];
@(posedge clk);
#1;data_in = testData5[615];
@(posedge clk);
#1;data_in = testData5[616];
@(posedge clk);
#1;data_in = testData5[617];
@(posedge clk);
#1;data_in = testData5[618];
@(posedge clk);
#1;data_in = testData5[619];
@(posedge clk);
#1;data_in = testData5[620];
@(posedge clk);
#1;data_in = testData5[621];
@(posedge clk);
#1;data_in = testData5[622];
@(posedge clk);
#1;data_in = testData5[623];
@(posedge clk);
#1;data_in = testData5[624];
@(posedge clk);
#1;data_in = testData5[625];
@(posedge clk);
#1;data_in = testData5[626];
@(posedge clk);
#1;data_in = testData5[627];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[628]; 
@(posedge clk);
#1;data_in = testData5[629];
@(posedge clk);
#1;data_in = testData5[630];
@(posedge clk);
#1;data_in = testData5[631];
@(posedge clk);
#1;data_in = testData5[632];
@(posedge clk);
#1;data_in = testData5[633];
@(posedge clk);
#1;data_in = testData5[634];
@(posedge clk);
#1;data_in = testData5[635];
@(posedge clk);
#1;data_in = testData5[636];
@(posedge clk);
#1;data_in = testData5[637];
@(posedge clk);
#1;data_in = testData5[638];
@(posedge clk);
#1;data_in = testData5[639];
@(posedge clk);
#1;data_in = testData5[640];
@(posedge clk);
#1;data_in = testData5[641];
@(posedge clk);
#1;data_in = testData5[642];
@(posedge clk);
#1;data_in = testData5[643];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[644]; 
@(posedge clk);
#1;data_in = testData5[645];
@(posedge clk);
#1;data_in = testData5[646];
@(posedge clk);
#1;data_in = testData5[647];
@(posedge clk);
#1;data_in = testData5[648];
@(posedge clk);
#1;data_in = testData5[649];
@(posedge clk);
#1;data_in = testData5[650];
@(posedge clk);
#1;data_in = testData5[651];
@(posedge clk);
#1;data_in = testData5[652];
@(posedge clk);
#1;data_in = testData5[653];
@(posedge clk);
#1;data_in = testData5[654];
@(posedge clk);
#1;data_in = testData5[655];
@(posedge clk);
#1;data_in = testData5[656];
@(posedge clk);
#1;data_in = testData5[657];
@(posedge clk);
#1;data_in = testData5[658];
@(posedge clk);
#1;data_in = testData5[659];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[660]; 
@(posedge clk);
#1;data_in = testData5[661];
@(posedge clk);
#1;data_in = testData5[662];
@(posedge clk);
#1;data_in = testData5[663];
@(posedge clk);
#1;data_in = testData5[664];
@(posedge clk);
#1;data_in = testData5[665];
@(posedge clk);
#1;data_in = testData5[666];
@(posedge clk);
#1;data_in = testData5[667];
@(posedge clk);
#1;data_in = testData5[668];
@(posedge clk);
#1;data_in = testData5[669];
@(posedge clk);
#1;data_in = testData5[670];
@(posedge clk);
#1;data_in = testData5[671];
@(posedge clk);
#1;data_in = testData5[672];
@(posedge clk);
#1;data_in = testData5[673];
@(posedge clk);
#1;data_in = testData5[674];
@(posedge clk);
#1;data_in = testData5[675];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[676]; 
@(posedge clk);
#1;data_in = testData5[677];
@(posedge clk);
#1;data_in = testData5[678];
@(posedge clk);
#1;data_in = testData5[679];
@(posedge clk);
#1;data_in = testData5[680];
@(posedge clk);
#1;data_in = testData5[681];
@(posedge clk);
#1;data_in = testData5[682];
@(posedge clk);
#1;data_in = testData5[683];
@(posedge clk);
#1;data_in = testData5[684];
@(posedge clk);
#1;data_in = testData5[685];
@(posedge clk);
#1;data_in = testData5[686];
@(posedge clk);
#1;data_in = testData5[687];
@(posedge clk);
#1;data_in = testData5[688];
@(posedge clk);
#1;data_in = testData5[689];
@(posedge clk);
#1;data_in = testData5[690];
@(posedge clk);
#1;data_in = testData5[691];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[692]; 
@(posedge clk);
#1;data_in = testData5[693];
@(posedge clk);
#1;data_in = testData5[694];
@(posedge clk);
#1;data_in = testData5[695];
@(posedge clk);
#1;data_in = testData5[696];
@(posedge clk);
#1;data_in = testData5[697];
@(posedge clk);
#1;data_in = testData5[698];
@(posedge clk);
#1;data_in = testData5[699];
@(posedge clk);
#1;data_in = testData5[700];
@(posedge clk);
#1;data_in = testData5[701];
@(posedge clk);
#1;data_in = testData5[702];
@(posedge clk);
#1;data_in = testData5[703];
@(posedge clk);
#1;data_in = testData5[704];
@(posedge clk);
#1;data_in = testData5[705];
@(posedge clk);
#1;data_in = testData5[706];
@(posedge clk);
#1;data_in = testData5[707];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[708]; 
@(posedge clk);
#1;data_in = testData5[709];
@(posedge clk);
#1;data_in = testData5[710];
@(posedge clk);
#1;data_in = testData5[711];
@(posedge clk);
#1;data_in = testData5[712];
@(posedge clk);
#1;data_in = testData5[713];
@(posedge clk);
#1;data_in = testData5[714];
@(posedge clk);
#1;data_in = testData5[715];
@(posedge clk);
#1;data_in = testData5[716];
@(posedge clk);
#1;data_in = testData5[717];
@(posedge clk);
#1;data_in = testData5[718];
@(posedge clk);
#1;data_in = testData5[719];
@(posedge clk);
#1;data_in = testData5[720];
@(posedge clk);
#1;data_in = testData5[721];
@(posedge clk);
#1;data_in = testData5[722];
@(posedge clk);
#1;data_in = testData5[723];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[724]; 
@(posedge clk);
#1;data_in = testData5[725];
@(posedge clk);
#1;data_in = testData5[726];
@(posedge clk);
#1;data_in = testData5[727];
@(posedge clk);
#1;data_in = testData5[728];
@(posedge clk);
#1;data_in = testData5[729];
@(posedge clk);
#1;data_in = testData5[730];
@(posedge clk);
#1;data_in = testData5[731];
@(posedge clk);
#1;data_in = testData5[732];
@(posedge clk);
#1;data_in = testData5[733];
@(posedge clk);
#1;data_in = testData5[734];
@(posedge clk);
#1;data_in = testData5[735];
@(posedge clk);
#1;data_in = testData5[736];
@(posedge clk);
#1;data_in = testData5[737];
@(posedge clk);
#1;data_in = testData5[738];
@(posedge clk);
#1;data_in = testData5[739];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[740]; 
@(posedge clk);
#1;data_in = testData5[741];
@(posedge clk);
#1;data_in = testData5[742];
@(posedge clk);
#1;data_in = testData5[743];
@(posedge clk);
#1;data_in = testData5[744];
@(posedge clk);
#1;data_in = testData5[745];
@(posedge clk);
#1;data_in = testData5[746];
@(posedge clk);
#1;data_in = testData5[747];
@(posedge clk);
#1;data_in = testData5[748];
@(posedge clk);
#1;data_in = testData5[749];
@(posedge clk);
#1;data_in = testData5[750];
@(posedge clk);
#1;data_in = testData5[751];
@(posedge clk);
#1;data_in = testData5[752];
@(posedge clk);
#1;data_in = testData5[753];
@(posedge clk);
#1;data_in = testData5[754];
@(posedge clk);
#1;data_in = testData5[755];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[756]; 
@(posedge clk);
#1;data_in = testData5[757];
@(posedge clk);
#1;data_in = testData5[758];
@(posedge clk);
#1;data_in = testData5[759];
@(posedge clk);
#1;data_in = testData5[760];
@(posedge clk);
#1;data_in = testData5[761];
@(posedge clk);
#1;data_in = testData5[762];
@(posedge clk);
#1;data_in = testData5[763];
@(posedge clk);
#1;data_in = testData5[764];
@(posedge clk);
#1;data_in = testData5[765];
@(posedge clk);
#1;data_in = testData5[766];
@(posedge clk);
#1;data_in = testData5[767];
@(posedge clk);
#1;data_in = testData5[768];
@(posedge clk);
#1;data_in = testData5[769];
@(posedge clk);
#1;data_in = testData5[770];
@(posedge clk);
#1;data_in = testData5[771];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[772]; 
@(posedge clk);
#1;data_in = testData5[773];
@(posedge clk);
#1;data_in = testData5[774];
@(posedge clk);
#1;data_in = testData5[775];
@(posedge clk);
#1;data_in = testData5[776];
@(posedge clk);
#1;data_in = testData5[777];
@(posedge clk);
#1;data_in = testData5[778];
@(posedge clk);
#1;data_in = testData5[779];
@(posedge clk);
#1;data_in = testData5[780];
@(posedge clk);
#1;data_in = testData5[781];
@(posedge clk);
#1;data_in = testData5[782];
@(posedge clk);
#1;data_in = testData5[783];
@(posedge clk);
#1;data_in = testData5[784];
@(posedge clk);
#1;data_in = testData5[785];
@(posedge clk);
#1;data_in = testData5[786];
@(posedge clk);
#1;data_in = testData5[787];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[788]; 
@(posedge clk);
#1;data_in = testData5[789];
@(posedge clk);
#1;data_in = testData5[790];
@(posedge clk);
#1;data_in = testData5[791];
@(posedge clk);
#1;data_in = testData5[792];
@(posedge clk);
#1;data_in = testData5[793];
@(posedge clk);
#1;data_in = testData5[794];
@(posedge clk);
#1;data_in = testData5[795];
@(posedge clk);
#1;data_in = testData5[796];
@(posedge clk);
#1;data_in = testData5[797];
@(posedge clk);
#1;data_in = testData5[798];
@(posedge clk);
#1;data_in = testData5[799];
@(posedge clk);
#1;data_in = testData5[800];
@(posedge clk);
#1;data_in = testData5[801];
@(posedge clk);
#1;data_in = testData5[802];
@(posedge clk);
#1;data_in = testData5[803];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
#1 ; loadMatrix =1;
@(posedge clk);
#1 ; loadMatrix =0;
data_in=testData5[804]; 
@(posedge clk);
#1;data_in = testData5[805];
@(posedge clk);
#1;data_in = testData5[806];
@(posedge clk);
#1;data_in = testData5[807];
@(posedge clk);
#1;data_in = testData5[808];
@(posedge clk);
#1;data_in = testData5[809];
@(posedge clk);
#1;data_in = testData5[810];
@(posedge clk);
#1;data_in = testData5[811];
@(posedge clk);
#1;data_in = testData5[812];
@(posedge clk);
#1;data_in = testData5[813];
@(posedge clk);
#1;data_in = testData5[814];
@(posedge clk);
#1;data_in = testData5[815];
@(posedge clk);
#1;data_in = testData5[816];
@(posedge clk);
#1;data_in = testData5[817];
@(posedge clk);
#1;data_in = testData5[818];
@(posedge clk);
#1;data_in = testData5[819];
@(posedge clk);
@(posedge clk);
#1; start=1;
@(posedge clk);
#1; start=0;
 
// wait for done signal and output  
@(posedge done);
 #1; qwerty=0;
@(posedge clk);
#1; $display("y[0] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[1] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[2] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
#1; $display("y[3] = %d" , data_out); $fdisplay(filehandle, "%d", data_out);
@(posedge clk);
$finish;
 end
 endmodule 
